LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY BasedVectorLFSR IS
	GENERIC ( n	: INTEGER	:= 2000			    -- number of bits
				);	 
	PORT (
		clk, rst, update	: IN STD_LOGIC; 
		dout				: OUT  STD_LOGIC_VECTOR (n-1 DOWNTO 0 )
	);
END ENTITY BasedVectorLFSR;

ARCHITECTURE behavioral OF BasedVectorLFSR IS

COMPONENT  regOne IS
	GENERIC (init : STD_LOGIC := '1');   -- initial value
	PORT (
		clk 				: IN  STD_LOGIC;
		regUpdate, regrst 	: IN  STD_LOGIC;
		din        			: IN  STD_LOGIC;
		dout        		: OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL interValIn : STD_LOGIC_VECTOR (n-1 DOWNTO 0);
SIGNAL interValOut : STD_LOGIC_VECTOR (n-1 DOWNTO 0);
SIGNAL interValOutR : STD_LOGIC_VECTOR (0 TO n-1);
CONSTANT congigSigniture : STD_LOGIC_VECTOR (n-1 DOWNTO 0) :=    "1000100001110111110011111110101101101111011010000101000100101101100101000000001011100000111111101001100011110110100111101011011100011010110101001110111000101101011111001101110001110001001011011001110110100100101101111010010011001101011000100011000011001000100111101010111111010110001001010011010111101110000010000001000010110100110100001101010101011101011010001100001101010100100001101000101110110000110001001110001100100010011111110000000011010001011010000000011101010010001110000111100110010110010000001111100000110111100011011110101011000001101000110111000111111001010011110011001111000110000011110011111001110010011100000110010011011010011100111100001000000010111011010000011110101010000000110111010011101011100001011101101011010110000010111011101000011001000011000000101100100001101111111100111001000010011101010101111001000100001111001011110101100000011010100011101100001001010011001011001101110100101100001011110010000000110011010001100010110011110111110010100100011000101010110111010100101011"; --"1010101011000011001011001000001001000110100100000010011011000001110101100010000001000111100011101100011001100110100010101100010001011111010110000011000010111011110110101000110101100100110110100001010010111100101010101000111011111101101111011111001111001010110000010110100001111110011100100000000110110110000000011011010111101011100110101100010100100011010011000001010111000000010001101101101011010110110011110000010000110110010110100011111001011110011010011101011010111100011001010111011111110101100110001110000011111111110110001011001111111110010101010010011101000011100111101011011000110101010101100000100001101010101000111111001001111101010000110001110110001010111000101100101010011110010101100010011011011111111100100111100010011100101010010000001100111011100101101011100010111001000110101111110111111010001000100101100011100010001011001100110111011010101010000010100000000101001000110011011011011100010011011001001011100000000000000001000010010101100101110110001001101010101101010001110000001100";

CONSTANT congigInitialvalues : STD_LOGIC_VECTOR (n-1 DOWNTO 0) := "0111011000100111101100100000001101100110010001101010010011010010111011001000000111000000111110100111100011000011001101110000110011011010100000001100001010000010100111111110100011010011111111111111011100101100101011111110011001000111101100001111001100101000111000100011100101110011111100101111000100000011100001001101010100001110101110110100101101100110101001001011011001111000011101010001110111000101111100010100111100110111110101000100110010100001011111111100010111011001010110001100001110011110000101000100100001000010000010010011011100111100100110100001100100010001111011101011000111101000100100011001111110100100010101010101110000010010000000100010111011011111011101101101111001000101111000110110011011111111110111010000000110111110000111100110001011000010110011111000111101011000010111101101001111011000010001100101110110001101100001110110110001000001001110011101110010100110011001011001010010101001111111000110110000101000111110110100010000110100010001000011010101000110001000111000010111001110";--"1111000000100110110100000110111010000101111100010011000110000110000100100100100010111110100100111000000001010111001001001000111010011010000001011010010100111000100010110111010111110010000101010100011101011111011100001011010100011100110110100001101100111100101111001001100100000011110111000110111000010001111100011110001110001010001011011011000000001010000001000001000011100010110011111101111000000010000111110001101011110111101010101010001110110110100100101011011011011110000111110110011000100110111010000011101100111010000010101011010111001011110110100000101100101111110011010011010010111000100100101100101101010001001110100010100001011100010111110010110011101000111110110001100100011100001110110000101111110011100100011011011101101110010101000101010100101011110011100100111100010011011100100101001010000110000101011100001110011111100011000011101010100001011010100101011110000100010001101001000000001011010001001001001000111010110101000010101011111110000010001010100111111100100011000110110101100110";

BEGIN

	regArr : FOR i IN 1 TO n-1 GENERATE
		Ireg : regOne 
			GENERIC map(congigInitialvalues(i))
			PORT map(clk,  update, rst, 
			interValIn(i), 	interValOut(i) 
					 );   
	END GENERATE regArr;
	xorchain : FOR i IN 1 TO n-1 GENERATE
	xorchain1: IF (congigSigniture(i) = '1') GENERATE
			interValIn(i) <= interValOut(i-1) XOR  interValOut(n-1);
		END GENERATE xorchain1;
	xorchain2: IF (congigSigniture(i) = '0') GENERATE
			interValIn(i) <= interValOut(i-1);
		END GENERATE xorchain2;
	END GENERATE xorchain;
	interValIn(0) <= interValOut(n-1);
	reg0 : regOne 
			GENERIC map(congigInitialvalues(0))
			PORT map(clk,  update, rst, 
			interValIn(0), 	interValOut(0) 
					 ); 
	--interValOutR <= interValOut;
	dout <= interValOut;--(0 TO n-1);

END ARCHITECTURE behavioral;