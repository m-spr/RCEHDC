LIBRARY IEEE; 
USE IEEE.STD_LOGIC_1164.ALL; 
USE IEEE.NUMERIC_STD.ALL; 
  
ENTITY connector IS 
	GENERIC(d : INTEGER := 1000; ----dimentionsize 
	p: INTEGER:= 1000 ); --- prunsize 
	PORT ( 
		input         : IN  STD_LOGIC_VECTOR (d-1 DOWNTO 0); 
		pruneoutput        : OUT  STD_LOGIC_VECTOR (p-1 DOWNTO 0)      
	);
END ENTITY connector;

ARCHITECTURE behavioral OF connector  IS
BEGIN
	 pruneoutput(335) <= input(992);
	 pruneoutput(334) <= input(991);
	 pruneoutput(333) <= input(984);
	 pruneoutput(332) <= input(981);
	 pruneoutput(331) <= input(980);
	 pruneoutput(330) <= input(979);
	 pruneoutput(329) <= input(973);
	 pruneoutput(328) <= input(970);
	 pruneoutput(327) <= input(969);
	 pruneoutput(326) <= input(965);
	 pruneoutput(325) <= input(964);
	 pruneoutput(324) <= input(963);
	 pruneoutput(323) <= input(959);
	 pruneoutput(322) <= input(958);
	 pruneoutput(321) <= input(954);
	 pruneoutput(320) <= input(953);
	 pruneoutput(319) <= input(952);
	 pruneoutput(318) <= input(951);
	 pruneoutput(317) <= input(943);
	 pruneoutput(316) <= input(942);
	 pruneoutput(315) <= input(941);
	 pruneoutput(314) <= input(937);
	 pruneoutput(313) <= input(936);
	 pruneoutput(312) <= input(929);
	 pruneoutput(311) <= input(928);
	 pruneoutput(310) <= input(927);
	 pruneoutput(309) <= input(926);
	 pruneoutput(308) <= input(925);
	 pruneoutput(307) <= input(924);
	 pruneoutput(306) <= input(923);
	 pruneoutput(305) <= input(893);
	 pruneoutput(304) <= input(886);
	 pruneoutput(303) <= input(885);
	 pruneoutput(302) <= input(884);
	 pruneoutput(301) <= input(883);
	 pruneoutput(300) <= input(882);
	 pruneoutput(299) <= input(880);
	 pruneoutput(298) <= input(879);
	 pruneoutput(297) <= input(877);
	 pruneoutput(296) <= input(869);
	 pruneoutput(295) <= input(868);
	 pruneoutput(294) <= input(865);
	 pruneoutput(293) <= input(862);
	 pruneoutput(292) <= input(857);
	 pruneoutput(291) <= input(856);
	 pruneoutput(290) <= input(855);
	 pruneoutput(289) <= input(854);
	 pruneoutput(288) <= input(852);
	 pruneoutput(287) <= input(851);
	 pruneoutput(286) <= input(850);
	 pruneoutput(285) <= input(848);
	 pruneoutput(284) <= input(847);
	 pruneoutput(283) <= input(846);
	 pruneoutput(282) <= input(845);
	 pruneoutput(281) <= input(839);
	 pruneoutput(280) <= input(837);
	 pruneoutput(279) <= input(832);
	 pruneoutput(278) <= input(831);
	 pruneoutput(277) <= input(830);
	 pruneoutput(276) <= input(825);
	 pruneoutput(275) <= input(824);
	 pruneoutput(274) <= input(820);
	 pruneoutput(273) <= input(819);
	 pruneoutput(272) <= input(818);
	 pruneoutput(271) <= input(817);
	 pruneoutput(270) <= input(813);
	 pruneoutput(269) <= input(810);
	 pruneoutput(268) <= input(807);
	 pruneoutput(267) <= input(802);
	 pruneoutput(266) <= input(801);
	 pruneoutput(265) <= input(800);
	 pruneoutput(264) <= input(798);
	 pruneoutput(263) <= input(797);
	 pruneoutput(262) <= input(784);
	 pruneoutput(261) <= input(783);
	 pruneoutput(260) <= input(782);
	 pruneoutput(259) <= input(781);
	 pruneoutput(258) <= input(769);
	 pruneoutput(257) <= input(768);
	 pruneoutput(256) <= input(742);
	 pruneoutput(255) <= input(741);
	 pruneoutput(254) <= input(740);
	 pruneoutput(253) <= input(734);
	 pruneoutput(252) <= input(733);
	 pruneoutput(251) <= input(732);
	 pruneoutput(250) <= input(731);
	 pruneoutput(249) <= input(730);
	 pruneoutput(248) <= input(721);
	 pruneoutput(247) <= input(713);
	 pruneoutput(246) <= input(712);
	 pruneoutput(245) <= input(705);
	 pruneoutput(244) <= input(704);
	 pruneoutput(243) <= input(703);
	 pruneoutput(242) <= input(701);
	 pruneoutput(241) <= input(696);
	 pruneoutput(240) <= input(695);
	 pruneoutput(239) <= input(694);
	 pruneoutput(238) <= input(693);
	 pruneoutput(237) <= input(677);
	 pruneoutput(236) <= input(669);
	 pruneoutput(235) <= input(668);
	 pruneoutput(234) <= input(661);
	 pruneoutput(233) <= input(660);
	 pruneoutput(232) <= input(657);
	 pruneoutput(231) <= input(656);
	 pruneoutput(230) <= input(655);
	 pruneoutput(229) <= input(654);
	 pruneoutput(228) <= input(649);
	 pruneoutput(227) <= input(648);
	 pruneoutput(226) <= input(647);
	 pruneoutput(225) <= input(642);
	 pruneoutput(224) <= input(641);
	 pruneoutput(223) <= input(640);
	 pruneoutput(222) <= input(639);
	 pruneoutput(221) <= input(638);
	 pruneoutput(220) <= input(637);
	 pruneoutput(219) <= input(636);
	 pruneoutput(218) <= input(635);
	 pruneoutput(217) <= input(634);
	 pruneoutput(216) <= input(633);
	 pruneoutput(215) <= input(628);
	 pruneoutput(214) <= input(627);
	 pruneoutput(213) <= input(626);
	 pruneoutput(212) <= input(622);
	 pruneoutput(211) <= input(621);
	 pruneoutput(210) <= input(620);
	 pruneoutput(209) <= input(619);
	 pruneoutput(208) <= input(617);
	 pruneoutput(207) <= input(608);
	 pruneoutput(206) <= input(603);
	 pruneoutput(205) <= input(602);
	 pruneoutput(204) <= input(601);
	 pruneoutput(203) <= input(600);
	 pruneoutput(202) <= input(599);
	 pruneoutput(201) <= input(597);
	 pruneoutput(200) <= input(596);
	 pruneoutput(199) <= input(595);
	 pruneoutput(198) <= input(594);
	 pruneoutput(197) <= input(589);
	 pruneoutput(196) <= input(588);
	 pruneoutput(195) <= input(587);
	 pruneoutput(194) <= input(586);
	 pruneoutput(193) <= input(585);
	 pruneoutput(192) <= input(583);
	 pruneoutput(191) <= input(582);
	 pruneoutput(190) <= input(574);
	 pruneoutput(189) <= input(573);
	 pruneoutput(188) <= input(568);
	 pruneoutput(187) <= input(554);
	 pruneoutput(186) <= input(553);
	 pruneoutput(185) <= input(552);
	 pruneoutput(184) <= input(551);
	 pruneoutput(183) <= input(550);
	 pruneoutput(182) <= input(549);
	 pruneoutput(181) <= input(531);
	 pruneoutput(180) <= input(530);
	 pruneoutput(179) <= input(529);
	 pruneoutput(178) <= input(528);
	 pruneoutput(177) <= input(527);
	 pruneoutput(176) <= input(526);
	 pruneoutput(175) <= input(525);
	 pruneoutput(174) <= input(523);
	 pruneoutput(173) <= input(522);
	 pruneoutput(172) <= input(521);
	 pruneoutput(171) <= input(520);
	 pruneoutput(170) <= input(519);
	 pruneoutput(169) <= input(518);
	 pruneoutput(168) <= input(516);
	 pruneoutput(167) <= input(515);
	 pruneoutput(166) <= input(477);
	 pruneoutput(165) <= input(476);
	 pruneoutput(164) <= input(469);
	 pruneoutput(163) <= input(462);
	 pruneoutput(162) <= input(455);
	 pruneoutput(161) <= input(445);
	 pruneoutput(160) <= input(438);
	 pruneoutput(159) <= input(437);
	 pruneoutput(158) <= input(435);
	 pruneoutput(157) <= input(429);
	 pruneoutput(156) <= input(428);
	 pruneoutput(155) <= input(426);
	 pruneoutput(154) <= input(425);
	 pruneoutput(153) <= input(422);
	 pruneoutput(152) <= input(414);
	 pruneoutput(151) <= input(409);
	 pruneoutput(150) <= input(407);
	 pruneoutput(149) <= input(404);
	 pruneoutput(148) <= input(403);
	 pruneoutput(147) <= input(396);
	 pruneoutput(146) <= input(390);
	 pruneoutput(145) <= input(389);
	 pruneoutput(144) <= input(388);
	 pruneoutput(143) <= input(381);
	 pruneoutput(142) <= input(380);
	 pruneoutput(141) <= input(379);
	 pruneoutput(140) <= input(378);
	 pruneoutput(139) <= input(377);
	 pruneoutput(138) <= input(373);
	 pruneoutput(137) <= input(372);
	 pruneoutput(136) <= input(371);
	 pruneoutput(135) <= input(370);
	 pruneoutput(134) <= input(367);
	 pruneoutput(133) <= input(360);
	 pruneoutput(132) <= input(359);
	 pruneoutput(131) <= input(358);
	 pruneoutput(130) <= input(351);
	 pruneoutput(129) <= input(349);
	 pruneoutput(128) <= input(348);
	 pruneoutput(127) <= input(347);
	 pruneoutput(126) <= input(333);
	 pruneoutput(125) <= input(332);
	 pruneoutput(124) <= input(331);
	 pruneoutput(123) <= input(330);
	 pruneoutput(122) <= input(321);
	 pruneoutput(121) <= input(316);
	 pruneoutput(120) <= input(315);
	 pruneoutput(119) <= input(314);
	 pruneoutput(118) <= input(313);
	 pruneoutput(117) <= input(303);
	 pruneoutput(116) <= input(302);
	 pruneoutput(115) <= input(299);
	 pruneoutput(114) <= input(298);
	 pruneoutput(113) <= input(294);
	 pruneoutput(112) <= input(293);
	 pruneoutput(111) <= input(292);
	 pruneoutput(110) <= input(291);
	 pruneoutput(109) <= input(284);
	 pruneoutput(108) <= input(283);
	 pruneoutput(107) <= input(282);
	 pruneoutput(106) <= input(272);
	 pruneoutput(105) <= input(271);
	 pruneoutput(104) <= input(267);
	 pruneoutput(103) <= input(266);
	 pruneoutput(102) <= input(264);
	 pruneoutput(101) <= input(263);
	 pruneoutput(100) <= input(262);
	 pruneoutput(99) <= input(261);
	 pruneoutput(98) <= input(260);
	 pruneoutput(97) <= input(259);
	 pruneoutput(96) <= input(258);
	 pruneoutput(95) <= input(256);
	 pruneoutput(94) <= input(250);
	 pruneoutput(93) <= input(249);
	 pruneoutput(92) <= input(233);
	 pruneoutput(91) <= input(232);
	 pruneoutput(90) <= input(231);
	 pruneoutput(89) <= input(230);
	 pruneoutput(88) <= input(229);
	 pruneoutput(87) <= input(228);
	 pruneoutput(86) <= input(227);
	 pruneoutput(85) <= input(226);
	 pruneoutput(84) <= input(225);
	 pruneoutput(83) <= input(222);
	 pruneoutput(82) <= input(221);
	 pruneoutput(81) <= input(211);
	 pruneoutput(80) <= input(206);
	 pruneoutput(79) <= input(205);
	 pruneoutput(78) <= input(204);
	 pruneoutput(77) <= input(202);
	 pruneoutput(76) <= input(199);
	 pruneoutput(75) <= input(198);
	 pruneoutput(74) <= input(191);
	 pruneoutput(73) <= input(190);
	 pruneoutput(72) <= input(187);
	 pruneoutput(71) <= input(185);
	 pruneoutput(70) <= input(184);
	 pruneoutput(69) <= input(181);
	 pruneoutput(68) <= input(180);
	 pruneoutput(67) <= input(179);
	 pruneoutput(66) <= input(176);
	 pruneoutput(65) <= input(175);
	 pruneoutput(64) <= input(174);
	 pruneoutput(63) <= input(163);
	 pruneoutput(62) <= input(151);
	 pruneoutput(61) <= input(150);
	 pruneoutput(60) <= input(149);
	 pruneoutput(59) <= input(141);
	 pruneoutput(58) <= input(138);
	 pruneoutput(57) <= input(137);
	 pruneoutput(56) <= input(136);
	 pruneoutput(55) <= input(135);
	 pruneoutput(54) <= input(134);
	 pruneoutput(53) <= input(133);
	 pruneoutput(52) <= input(127);
	 pruneoutput(51) <= input(126);
	 pruneoutput(50) <= input(125);
	 pruneoutput(49) <= input(124);
	 pruneoutput(48) <= input(123);
	 pruneoutput(47) <= input(113);
	 pruneoutput(46) <= input(112);
	 pruneoutput(45) <= input(111);
	 pruneoutput(44) <= input(110);
	 pruneoutput(43) <= input(109);
	 pruneoutput(42) <= input(104);
	 pruneoutput(41) <= input(100);
	 pruneoutput(40) <= input(97);
	 pruneoutput(39) <= input(96);
	 pruneoutput(38) <= input(95);
	 pruneoutput(37) <= input(94);
	 pruneoutput(36) <= input(93);
	 pruneoutput(35) <= input(86);
	 pruneoutput(34) <= input(83);
	 pruneoutput(33) <= input(78);
	 pruneoutput(32) <= input(77);
	 pruneoutput(31) <= input(76);
	 pruneoutput(30) <= input(70);
	 pruneoutput(29) <= input(69);
	 pruneoutput(28) <= input(68);
	 pruneoutput(27) <= input(67);
	 pruneoutput(26) <= input(66);
	 pruneoutput(25) <= input(63);
	 pruneoutput(24) <= input(62);
	 pruneoutput(23) <= input(61);
	 pruneoutput(22) <= input(60);
	 pruneoutput(21) <= input(47);
	 pruneoutput(20) <= input(46);
	 pruneoutput(19) <= input(40);
	 pruneoutput(18) <= input(36);
	 pruneoutput(17) <= input(35);
	 pruneoutput(16) <= input(29);
	 pruneoutput(15) <= input(28);
	 pruneoutput(14) <= input(26);
	 pruneoutput(13) <= input(25);
	 pruneoutput(12) <= input(23);
	 pruneoutput(11) <= input(22);
	 pruneoutput(10) <= input(21);
	 pruneoutput(9) <= input(18);
	 pruneoutput(8) <= input(17);
	 pruneoutput(7) <= input(15);
	 pruneoutput(6) <= input(14);
	 pruneoutput(5) <= input(13);
	 pruneoutput(4) <= input(11);
	 pruneoutput(3) <= input(10);
	 pruneoutput(2) <= input(8);
	 pruneoutput(1) <= input(4);
	 pruneoutput(0) <= input(3);

END ARCHITECTURE behavioral;