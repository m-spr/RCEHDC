LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY BasedVectorLFSR IS
	GENERIC ( n	: INTEGER	:= 2000			    -- number of bits
				);	 
	PORT (
		clk, rst, update	: IN STD_LOGIC; 
		congigSignitureIn , congigInitialvaluesIn : IN STD_LOGIC_VECTOR (n-1 DOWNTO 0 );
		dout				: OUT  STD_LOGIC_VECTOR (n-1 DOWNTO 0 )
	);
END ENTITY BasedVectorLFSR;

ARCHITECTURE behavioral OF BasedVectorLFSR IS

COMPONENT  regOne IS
	GENERIC (init : STD_LOGIC := '1');   -- initial value
	PORT (
		clk 				: IN  STD_LOGIC;
		regUpdate, regrst 	: IN  STD_LOGIC;
		din        			: IN  STD_LOGIC;
		dout        		: OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL interValIn : STD_LOGIC_VECTOR (n-1 DOWNTO 0);
SIGNAL interValOut : STD_LOGIC_VECTOR (n-1 DOWNTO 0);
SIGNAL interValOutR : STD_LOGIC_VECTOR (0 TO n-1);
CONSTANT congigSigniture : STD_LOGIC_VECTOR (n-1 DOWNTO 0) :=    "10100101110100010011010111001101110110100110000100110101011101010010001010100110111100001110000111001001001101101010000100011110110001011000001001100000111111100011110001110110111110101001001000110111001001101001110001000010100111001111010111001101101111111000101110110100101101111011110101001111111110000100010100110010111000111110011110001000010111011100101101001011101101111101010111001011001110110110101100001001110001001111001000100110000010110111110000100100111011000011110100001111010110111011011111100011011100110101000100110000011111001111001110111010101000111111111101111000101110010111100111000001010010100010000100011011101111011111101011011101110000110111001001111010111001001010001101110101011100001100000101100110011101011111111100100100011100111001011011011000000110111011011000100010010110000101101111100111100001101111001001011101100001000001011110000101001001011010100101100001101110100000001001011111010111110010111111011110101110010101100111010001010101110110000001010100001101001001000111001001110110000010001000111000000110001110101110111010010011000100110010110011000110101011"; --"1010101011000011001011001000001001000110100100000010011011000001110101100010000001000111100011101100011001100110100010101100010001011111010110000011000010111011110110101000110101100100110110100001010010111100101010101000111011111101101111011111001111001010110000010110100001111110011100100000000110110110000000011011010111101011100110101100010100100011010011000001010111000000010001101101101011010110110011110000010000110110010110100011111001011110011010011101011010111100011001010111011111110101100110001110000011111111110110001011001111111110010101010010011101000011100111101011011000110101010101100000100001101010101000111111001001111101010000110001110110001010111000101100101010011110010101100010011011011111111100100111100010011100101010010000001100111011100101101011100010111001000110101111110111111010001000100101100011100010001011001100110111011010101010000010100000000101001000110011011011011100010011011001001011100000000000000001000010010101100101110110001001101010101101010001110000001100";

CONSTANT congigInitialvalues : STD_LOGIC_VECTOR (n-1 DOWNTO 0) := "01100011101011100011100001000100011111001011101100110011111000101000110110111011111101000000101101111010101111111000110001110100011101010110100010001010111110101101011010000001011111111001101010001101011001001100101001110010101000101111000110000001010011001110001000100000100010110100111010100000011001101011111101010110000111100110011001110110110010101101000001101010001110101101011011110111111010000100001010100000110010111101000100101111110111010111001011111001000111011001111101010010000010110101100101000101000101001010101110110100101000111111110011111110110000110111000101001011110010101011111100111001011010100100000001100100000000100011111010101011001111011010111000011000001001011101000010001111110001101001111001111100010010111001000001101011001101011011100111000101011111111011111110010001000111001100000011001101111100001101001000101100101100010011000001100101011010101101010110011010011100101101100111100010101101101111101000101000111011011001000000000111100001101100001011001110001010000111111110001111111101100010001101100000110100001111010001110110000101010000000100010001011100110100";--"1111000000100110110100000110111010000101111100010011000110000110000100100100100010111110100100111000000001010111001001001000111010011010000001011010010100111000100010110111010111110010000101010100011101011111011100001011010100011100110110100001101100111100101111001001100100000011110111000110111000010001111100011110001110001010001011011011000000001010000001000001000011100010110011111101111000000010000111110001101011110111101010101010001110110110100100101011011011011110000111110110011000100110111010000011101100111010000010101011010111001011110110100000101100101111110011010011010010111000100100101100101101010001001110100010100001011100010111110010110011101000111110110001100100011100001110110000101111110011100100011011011101101110010101000101010100101011110011100100111100010011011100100101001010000110000101011100001110011111100011000011101010100001011010100101011110000100010001101001000000001011010001001001001000111010110101000010101011111110000010001010100111111100100011000110110101100110";

BEGIN

	regArr : FOR i IN 1 TO n-1 GENERATE
		Ireg : regOne 
			GENERIC map(congigInitialvalues(i))
			PORT map(clk,  update, rst, 
			interValIn(i), 	interValOut(i) 
					 );   
	END GENERATE regArr;
	xorchain : FOR i IN 1 TO n-1 GENERATE
	xorchain1: IF (congigSigniture(i) = '1') GENERATE
			interValIn(i) <= interValOut(i-1) XOR  interValOut(n-1);
		END GENERATE xorchain1;
	xorchain2: IF (congigSigniture(i) = '0') GENERATE
			interValIn(i) <= interValOut(i-1);
		END GENERATE xorchain2;
	END GENERATE xorchain;
	interValIn(0) <= interValOut(n-1);
	reg0 : regOne 
			GENERIC map(congigInitialvalues(0))
			PORT map(clk,  update, rst, 
			interValIn(0), 	interValOut(0) 
					 ); 
	--interValOutR <= interValOut;
	dout <= interValOut;--(0 TO n-1);

END ARCHITECTURE behavioral;