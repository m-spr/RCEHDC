LIBRARY IEEE; 
USE IEEE.STD_LOGIC_1164.ALL; 
USE IEEE.NUMERIC_STD.ALL; 
  
ENTITY connector IS 
	GENERIC(d : INTEGER := 1000; ----dimentionsize 
	p: INTEGER:= 1000 ); --- prunsize 
	PORT ( 
		input         : IN  STD_LOGIC_VECTOR (d-1 DOWNTO 0); 
		pruneoutput        : OUT  STD_LOGIC_VECTOR (p-1 DOWNTO 0)      
	);
END ENTITY connector;

ARCHITECTURE behavioral OF connector  IS
BEGIN
	 pruneoutput(386) <= input(999);
	 pruneoutput(385) <= input(997);
	 pruneoutput(384) <= input(996);
	 pruneoutput(383) <= input(980);
	 pruneoutput(382) <= input(979);
	 pruneoutput(381) <= input(978);
	 pruneoutput(380) <= input(977);
	 pruneoutput(379) <= input(971);
	 pruneoutput(378) <= input(970);
	 pruneoutput(377) <= input(968);
	 pruneoutput(376) <= input(967);
	 pruneoutput(375) <= input(956);
	 pruneoutput(374) <= input(943);
	 pruneoutput(373) <= input(938);
	 pruneoutput(372) <= input(937);
	 pruneoutput(371) <= input(936);
	 pruneoutput(370) <= input(926);
	 pruneoutput(369) <= input(925);
	 pruneoutput(368) <= input(915);
	 pruneoutput(367) <= input(914);
	 pruneoutput(366) <= input(912);
	 pruneoutput(365) <= input(911);
	 pruneoutput(364) <= input(910);
	 pruneoutput(363) <= input(904);
	 pruneoutput(362) <= input(903);
	 pruneoutput(361) <= input(902);
	 pruneoutput(360) <= input(898);
	 pruneoutput(359) <= input(894);
	 pruneoutput(358) <= input(893);
	 pruneoutput(357) <= input(892);
	 pruneoutput(356) <= input(891);
	 pruneoutput(355) <= input(890);
	 pruneoutput(354) <= input(889);
	 pruneoutput(353) <= input(888);
	 pruneoutput(352) <= input(887);
	 pruneoutput(351) <= input(886);
	 pruneoutput(350) <= input(885);
	 pruneoutput(349) <= input(884);
	 pruneoutput(348) <= input(882);
	 pruneoutput(347) <= input(873);
	 pruneoutput(346) <= input(870);
	 pruneoutput(345) <= input(867);
	 pruneoutput(344) <= input(866);
	 pruneoutput(343) <= input(865);
	 pruneoutput(342) <= input(858);
	 pruneoutput(341) <= input(857);
	 pruneoutput(340) <= input(856);
	 pruneoutput(339) <= input(855);
	 pruneoutput(338) <= input(854);
	 pruneoutput(337) <= input(851);
	 pruneoutput(336) <= input(838);
	 pruneoutput(335) <= input(837);
	 pruneoutput(334) <= input(836);
	 pruneoutput(333) <= input(835);
	 pruneoutput(332) <= input(833);
	 pruneoutput(331) <= input(832);
	 pruneoutput(330) <= input(831);
	 pruneoutput(329) <= input(830);
	 pruneoutput(328) <= input(829);
	 pruneoutput(327) <= input(828);
	 pruneoutput(326) <= input(827);
	 pruneoutput(325) <= input(826);
	 pruneoutput(324) <= input(820);
	 pruneoutput(323) <= input(818);
	 pruneoutput(322) <= input(810);
	 pruneoutput(321) <= input(809);
	 pruneoutput(320) <= input(808);
	 pruneoutput(319) <= input(807);
	 pruneoutput(318) <= input(806);
	 pruneoutput(317) <= input(805);
	 pruneoutput(316) <= input(803);
	 pruneoutput(315) <= input(802);
	 pruneoutput(314) <= input(793);
	 pruneoutput(313) <= input(792);
	 pruneoutput(312) <= input(791);
	 pruneoutput(311) <= input(789);
	 pruneoutput(310) <= input(788);
	 pruneoutput(309) <= input(785);
	 pruneoutput(308) <= input(779);
	 pruneoutput(307) <= input(777);
	 pruneoutput(306) <= input(775);
	 pruneoutput(305) <= input(772);
	 pruneoutput(304) <= input(771);
	 pruneoutput(303) <= input(770);
	 pruneoutput(302) <= input(768);
	 pruneoutput(301) <= input(756);
	 pruneoutput(300) <= input(755);
	 pruneoutput(299) <= input(754);
	 pruneoutput(298) <= input(753);
	 pruneoutput(297) <= input(752);
	 pruneoutput(296) <= input(746);
	 pruneoutput(295) <= input(745);
	 pruneoutput(294) <= input(744);
	 pruneoutput(293) <= input(743);
	 pruneoutput(292) <= input(732);
	 pruneoutput(291) <= input(731);
	 pruneoutput(290) <= input(722);
	 pruneoutput(289) <= input(721);
	 pruneoutput(288) <= input(720);
	 pruneoutput(287) <= input(710);
	 pruneoutput(286) <= input(702);
	 pruneoutput(285) <= input(701);
	 pruneoutput(284) <= input(700);
	 pruneoutput(283) <= input(699);
	 pruneoutput(282) <= input(698);
	 pruneoutput(281) <= input(697);
	 pruneoutput(280) <= input(696);
	 pruneoutput(279) <= input(695);
	 pruneoutput(278) <= input(694);
	 pruneoutput(277) <= input(692);
	 pruneoutput(276) <= input(691);
	 pruneoutput(275) <= input(690);
	 pruneoutput(274) <= input(676);
	 pruneoutput(273) <= input(675);
	 pruneoutput(272) <= input(674);
	 pruneoutput(271) <= input(673);
	 pruneoutput(270) <= input(671);
	 pruneoutput(269) <= input(670);
	 pruneoutput(268) <= input(669);
	 pruneoutput(267) <= input(665);
	 pruneoutput(266) <= input(664);
	 pruneoutput(265) <= input(656);
	 pruneoutput(264) <= input(655);
	 pruneoutput(263) <= input(654);
	 pruneoutput(262) <= input(653);
	 pruneoutput(261) <= input(650);
	 pruneoutput(260) <= input(649);
	 pruneoutput(259) <= input(648);
	 pruneoutput(258) <= input(640);
	 pruneoutput(257) <= input(639);
	 pruneoutput(256) <= input(634);
	 pruneoutput(255) <= input(632);
	 pruneoutput(254) <= input(631);
	 pruneoutput(253) <= input(630);
	 pruneoutput(252) <= input(628);
	 pruneoutput(251) <= input(627);
	 pruneoutput(250) <= input(626);
	 pruneoutput(249) <= input(625);
	 pruneoutput(248) <= input(624);
	 pruneoutput(247) <= input(623);
	 pruneoutput(246) <= input(622);
	 pruneoutput(245) <= input(621);
	 pruneoutput(244) <= input(620);
	 pruneoutput(243) <= input(619);
	 pruneoutput(242) <= input(618);
	 pruneoutput(241) <= input(617);
	 pruneoutput(240) <= input(616);
	 pruneoutput(239) <= input(615);
	 pruneoutput(238) <= input(603);
	 pruneoutput(237) <= input(600);
	 pruneoutput(236) <= input(595);
	 pruneoutput(235) <= input(594);
	 pruneoutput(234) <= input(587);
	 pruneoutput(233) <= input(584);
	 pruneoutput(232) <= input(583);
	 pruneoutput(231) <= input(577);
	 pruneoutput(230) <= input(575);
	 pruneoutput(229) <= input(574);
	 pruneoutput(228) <= input(573);
	 pruneoutput(227) <= input(572);
	 pruneoutput(226) <= input(571);
	 pruneoutput(225) <= input(570);
	 pruneoutput(224) <= input(569);
	 pruneoutput(223) <= input(568);
	 pruneoutput(222) <= input(567);
	 pruneoutput(221) <= input(566);
	 pruneoutput(220) <= input(565);
	 pruneoutput(219) <= input(564);
	 pruneoutput(218) <= input(563);
	 pruneoutput(217) <= input(561);
	 pruneoutput(216) <= input(560);
	 pruneoutput(215) <= input(558);
	 pruneoutput(214) <= input(555);
	 pruneoutput(213) <= input(554);
	 pruneoutput(212) <= input(539);
	 pruneoutput(211) <= input(538);
	 pruneoutput(210) <= input(537);
	 pruneoutput(209) <= input(535);
	 pruneoutput(208) <= input(534);
	 pruneoutput(207) <= input(533);
	 pruneoutput(206) <= input(532);
	 pruneoutput(205) <= input(531);
	 pruneoutput(204) <= input(516);
	 pruneoutput(203) <= input(515);
	 pruneoutput(202) <= input(514);
	 pruneoutput(201) <= input(513);
	 pruneoutput(200) <= input(505);
	 pruneoutput(199) <= input(500);
	 pruneoutput(198) <= input(499);
	 pruneoutput(197) <= input(497);
	 pruneoutput(196) <= input(482);
	 pruneoutput(195) <= input(481);
	 pruneoutput(194) <= input(480);
	 pruneoutput(193) <= input(472);
	 pruneoutput(192) <= input(471);
	 pruneoutput(191) <= input(467);
	 pruneoutput(190) <= input(466);
	 pruneoutput(189) <= input(465);
	 pruneoutput(188) <= input(464);
	 pruneoutput(187) <= input(463);
	 pruneoutput(186) <= input(448);
	 pruneoutput(185) <= input(447);
	 pruneoutput(184) <= input(444);
	 pruneoutput(183) <= input(443);
	 pruneoutput(182) <= input(442);
	 pruneoutput(181) <= input(432);
	 pruneoutput(180) <= input(431);
	 pruneoutput(179) <= input(430);
	 pruneoutput(178) <= input(428);
	 pruneoutput(177) <= input(424);
	 pruneoutput(176) <= input(420);
	 pruneoutput(175) <= input(413);
	 pruneoutput(174) <= input(412);
	 pruneoutput(173) <= input(411);
	 pruneoutput(172) <= input(410);
	 pruneoutput(171) <= input(407);
	 pruneoutput(170) <= input(406);
	 pruneoutput(169) <= input(405);
	 pruneoutput(168) <= input(404);
	 pruneoutput(167) <= input(403);
	 pruneoutput(166) <= input(402);
	 pruneoutput(165) <= input(401);
	 pruneoutput(164) <= input(400);
	 pruneoutput(163) <= input(399);
	 pruneoutput(162) <= input(398);
	 pruneoutput(161) <= input(396);
	 pruneoutput(160) <= input(395);
	 pruneoutput(159) <= input(391);
	 pruneoutput(158) <= input(390);
	 pruneoutput(157) <= input(388);
	 pruneoutput(156) <= input(387);
	 pruneoutput(155) <= input(386);
	 pruneoutput(154) <= input(385);
	 pruneoutput(153) <= input(375);
	 pruneoutput(152) <= input(369);
	 pruneoutput(151) <= input(367);
	 pruneoutput(150) <= input(350);
	 pruneoutput(149) <= input(349);
	 pruneoutput(148) <= input(348);
	 pruneoutput(147) <= input(346);
	 pruneoutput(146) <= input(334);
	 pruneoutput(145) <= input(331);
	 pruneoutput(144) <= input(330);
	 pruneoutput(143) <= input(327);
	 pruneoutput(142) <= input(326);
	 pruneoutput(141) <= input(324);
	 pruneoutput(140) <= input(323);
	 pruneoutput(139) <= input(322);
	 pruneoutput(138) <= input(320);
	 pruneoutput(137) <= input(310);
	 pruneoutput(136) <= input(309);
	 pruneoutput(135) <= input(298);
	 pruneoutput(134) <= input(297);
	 pruneoutput(133) <= input(295);
	 pruneoutput(132) <= input(294);
	 pruneoutput(131) <= input(293);
	 pruneoutput(130) <= input(292);
	 pruneoutput(129) <= input(291);
	 pruneoutput(128) <= input(290);
	 pruneoutput(127) <= input(289);
	 pruneoutput(126) <= input(288);
	 pruneoutput(125) <= input(287);
	 pruneoutput(124) <= input(286);
	 pruneoutput(123) <= input(285);
	 pruneoutput(122) <= input(284);
	 pruneoutput(121) <= input(283);
	 pruneoutput(120) <= input(282);
	 pruneoutput(119) <= input(281);
	 pruneoutput(118) <= input(278);
	 pruneoutput(117) <= input(277);
	 pruneoutput(116) <= input(276);
	 pruneoutput(115) <= input(275);
	 pruneoutput(114) <= input(274);
	 pruneoutput(113) <= input(268);
	 pruneoutput(112) <= input(267);
	 pruneoutput(111) <= input(266);
	 pruneoutput(110) <= input(265);
	 pruneoutput(109) <= input(263);
	 pruneoutput(108) <= input(262);
	 pruneoutput(107) <= input(261);
	 pruneoutput(106) <= input(260);
	 pruneoutput(105) <= input(259);
	 pruneoutput(104) <= input(258);
	 pruneoutput(103) <= input(244);
	 pruneoutput(102) <= input(243);
	 pruneoutput(101) <= input(242);
	 pruneoutput(100) <= input(240);
	 pruneoutput(99) <= input(234);
	 pruneoutput(98) <= input(233);
	 pruneoutput(97) <= input(231);
	 pruneoutput(96) <= input(230);
	 pruneoutput(95) <= input(229);
	 pruneoutput(94) <= input(228);
	 pruneoutput(93) <= input(227);
	 pruneoutput(92) <= input(225);
	 pruneoutput(91) <= input(218);
	 pruneoutput(90) <= input(217);
	 pruneoutput(89) <= input(216);
	 pruneoutput(88) <= input(213);
	 pruneoutput(87) <= input(212);
	 pruneoutput(86) <= input(211);
	 pruneoutput(85) <= input(210);
	 pruneoutput(84) <= input(209);
	 pruneoutput(83) <= input(208);
	 pruneoutput(82) <= input(207);
	 pruneoutput(81) <= input(206);
	 pruneoutput(80) <= input(205);
	 pruneoutput(79) <= input(204);
	 pruneoutput(78) <= input(198);
	 pruneoutput(77) <= input(191);
	 pruneoutput(76) <= input(190);
	 pruneoutput(75) <= input(187);
	 pruneoutput(74) <= input(184);
	 pruneoutput(73) <= input(171);
	 pruneoutput(72) <= input(170);
	 pruneoutput(71) <= input(169);
	 pruneoutput(70) <= input(162);
	 pruneoutput(69) <= input(155);
	 pruneoutput(68) <= input(154);
	 pruneoutput(67) <= input(152);
	 pruneoutput(66) <= input(151);
	 pruneoutput(65) <= input(150);
	 pruneoutput(64) <= input(149);
	 pruneoutput(63) <= input(148);
	 pruneoutput(62) <= input(146);
	 pruneoutput(61) <= input(145);
	 pruneoutput(60) <= input(142);
	 pruneoutput(59) <= input(139);
	 pruneoutput(58) <= input(134);
	 pruneoutput(57) <= input(132);
	 pruneoutput(56) <= input(131);
	 pruneoutput(55) <= input(128);
	 pruneoutput(54) <= input(127);
	 pruneoutput(53) <= input(126);
	 pruneoutput(52) <= input(116);
	 pruneoutput(51) <= input(115);
	 pruneoutput(50) <= input(108);
	 pruneoutput(49) <= input(107);
	 pruneoutput(48) <= input(102);
	 pruneoutput(47) <= input(101);
	 pruneoutput(46) <= input(100);
	 pruneoutput(45) <= input(99);
	 pruneoutput(44) <= input(98);
	 pruneoutput(43) <= input(97);
	 pruneoutput(42) <= input(93);
	 pruneoutput(41) <= input(87);
	 pruneoutput(40) <= input(86);
	 pruneoutput(39) <= input(85);
	 pruneoutput(38) <= input(84);
	 pruneoutput(37) <= input(83);
	 pruneoutput(36) <= input(82);
	 pruneoutput(35) <= input(75);
	 pruneoutput(34) <= input(69);
	 pruneoutput(33) <= input(68);
	 pruneoutput(32) <= input(65);
	 pruneoutput(31) <= input(64);
	 pruneoutput(30) <= input(62);
	 pruneoutput(29) <= input(61);
	 pruneoutput(28) <= input(60);
	 pruneoutput(27) <= input(59);
	 pruneoutput(26) <= input(58);
	 pruneoutput(25) <= input(57);
	 pruneoutput(24) <= input(56);
	 pruneoutput(23) <= input(55);
	 pruneoutput(22) <= input(54);
	 pruneoutput(21) <= input(53);
	 pruneoutput(20) <= input(49);
	 pruneoutput(19) <= input(48);
	 pruneoutput(18) <= input(47);
	 pruneoutput(17) <= input(41);
	 pruneoutput(16) <= input(32);
	 pruneoutput(15) <= input(24);
	 pruneoutput(14) <= input(23);
	 pruneoutput(13) <= input(22);
	 pruneoutput(12) <= input(21);
	 pruneoutput(11) <= input(17);
	 pruneoutput(10) <= input(16);
	 pruneoutput(9) <= input(14);
	 pruneoutput(8) <= input(13);
	 pruneoutput(7) <= input(12);
	 pruneoutput(6) <= input(10);
	 pruneoutput(5) <= input(9);
	 pruneoutput(4) <= input(8);
	 pruneoutput(3) <= input(6);
	 pruneoutput(2) <= input(5);
	 pruneoutput(1) <= input(4);
	 pruneoutput(0) <= input(0);

END ARCHITECTURE behavioral;