LIBRARY IEEE; 
USE IEEE.STD_LOGIC_1164.ALL; 
USE IEEE.NUMERIC_STD.ALL; 
  
ENTITY connector IS 
	PORT ( 
		input         : IN  STD_LOGIC_VECTOR (999 DOWNTO 0); 
		pruneoutput        : OUT  STD_LOGIC_VECTOR (645 DOWNTO 0)      
	);
END ENTITY connector;

ARCHITECTURE behavioral OF connector  IS
BEGIN
pruneoutput(0) <= input(0);
pruneoutput(1) <= input(1);
pruneoutput(2) <= input(2);
pruneoutput(3) <= input(4);
pruneoutput(4) <= input(5);
pruneoutput(5) <= input(6);
pruneoutput(6) <= input(13);
pruneoutput(7) <= input(14);
pruneoutput(8) <= input(15);
pruneoutput(9) <= input(18);
pruneoutput(10) <= input(19);
pruneoutput(11) <= input(20);
pruneoutput(12) <= input(21);
pruneoutput(13) <= input(22);
pruneoutput(14) <= input(23);
pruneoutput(15) <= input(25);
pruneoutput(16) <= input(26);
pruneoutput(17) <= input(27);
pruneoutput(18) <= input(28);
pruneoutput(19) <= input(29);
pruneoutput(20) <= input(33);
pruneoutput(21) <= input(35);
pruneoutput(22) <= input(37);
pruneoutput(23) <= input(39);
pruneoutput(24) <= input(40);
pruneoutput(25) <= input(41);
pruneoutput(26) <= input(42);
pruneoutput(27) <= input(43);
pruneoutput(28) <= input(44);
pruneoutput(29) <= input(48);
pruneoutput(30) <= input(49);
pruneoutput(31) <= input(52);
pruneoutput(32) <= input(56);
pruneoutput(33) <= input(57);
pruneoutput(34) <= input(58);
pruneoutput(35) <= input(59);
pruneoutput(36) <= input(60);
pruneoutput(37) <= input(63);
pruneoutput(38) <= input(64);
pruneoutput(39) <= input(65);
pruneoutput(40) <= input(66);
pruneoutput(41) <= input(67);
pruneoutput(42) <= input(68);
pruneoutput(43) <= input(69);
pruneoutput(44) <= input(73);
pruneoutput(45) <= input(74);
pruneoutput(46) <= input(75);
pruneoutput(47) <= input(76);
pruneoutput(48) <= input(77);
pruneoutput(49) <= input(78);
pruneoutput(50) <= input(80);
pruneoutput(51) <= input(81);
pruneoutput(52) <= input(82);
pruneoutput(53) <= input(83);
pruneoutput(54) <= input(84);
pruneoutput(55) <= input(85);
pruneoutput(56) <= input(86);
pruneoutput(57) <= input(87);
pruneoutput(58) <= input(88);
pruneoutput(59) <= input(89);
pruneoutput(60) <= input(91);
pruneoutput(61) <= input(92);
pruneoutput(62) <= input(93);
pruneoutput(63) <= input(94);
pruneoutput(64) <= input(95);
pruneoutput(65) <= input(103);
pruneoutput(66) <= input(104);
pruneoutput(67) <= input(105);
pruneoutput(68) <= input(106);
pruneoutput(69) <= input(108);
pruneoutput(70) <= input(109);
pruneoutput(71) <= input(110);
pruneoutput(72) <= input(112);
pruneoutput(73) <= input(113);
pruneoutput(74) <= input(114);
pruneoutput(75) <= input(115);
pruneoutput(76) <= input(116);
pruneoutput(77) <= input(118);
pruneoutput(78) <= input(121);
pruneoutput(79) <= input(122);
pruneoutput(80) <= input(127);
pruneoutput(81) <= input(128);
pruneoutput(82) <= input(129);
pruneoutput(83) <= input(133);
pruneoutput(84) <= input(134);
pruneoutput(85) <= input(135);
pruneoutput(86) <= input(136);
pruneoutput(87) <= input(137);
pruneoutput(88) <= input(138);
pruneoutput(89) <= input(141);
pruneoutput(90) <= input(146);
pruneoutput(91) <= input(147);
pruneoutput(92) <= input(148);
pruneoutput(93) <= input(149);
pruneoutput(94) <= input(150);
pruneoutput(95) <= input(151);
pruneoutput(96) <= input(152);
pruneoutput(97) <= input(154);
pruneoutput(98) <= input(155);
pruneoutput(99) <= input(156);
pruneoutput(100) <= input(157);
pruneoutput(101) <= input(158);
pruneoutput(102) <= input(159);
pruneoutput(103) <= input(160);
pruneoutput(104) <= input(161);
pruneoutput(105) <= input(165);
pruneoutput(106) <= input(171);
pruneoutput(107) <= input(172);
pruneoutput(108) <= input(173);
pruneoutput(109) <= input(179);
pruneoutput(110) <= input(181);
pruneoutput(111) <= input(184);
pruneoutput(112) <= input(185);
pruneoutput(113) <= input(186);
pruneoutput(114) <= input(187);
pruneoutput(115) <= input(191);
pruneoutput(116) <= input(192);
pruneoutput(117) <= input(193);
pruneoutput(118) <= input(196);
pruneoutput(119) <= input(199);
pruneoutput(120) <= input(200);
pruneoutput(121) <= input(203);
pruneoutput(122) <= input(204);
pruneoutput(123) <= input(206);
pruneoutput(124) <= input(207);
pruneoutput(125) <= input(210);
pruneoutput(126) <= input(211);
pruneoutput(127) <= input(217);
pruneoutput(128) <= input(218);
pruneoutput(129) <= input(219);
pruneoutput(130) <= input(220);
pruneoutput(131) <= input(225);
pruneoutput(132) <= input(228);
pruneoutput(133) <= input(229);
pruneoutput(134) <= input(230);
pruneoutput(135) <= input(231);
pruneoutput(136) <= input(232);
pruneoutput(137) <= input(233);
pruneoutput(138) <= input(234);
pruneoutput(139) <= input(235);
pruneoutput(140) <= input(236);
pruneoutput(141) <= input(237);
pruneoutput(142) <= input(239);
pruneoutput(143) <= input(240);
pruneoutput(144) <= input(241);
pruneoutput(145) <= input(242);
pruneoutput(146) <= input(243);
pruneoutput(147) <= input(244);
pruneoutput(148) <= input(245);
pruneoutput(149) <= input(249);
pruneoutput(150) <= input(250);
pruneoutput(151) <= input(253);
pruneoutput(152) <= input(254);
pruneoutput(153) <= input(261);
pruneoutput(154) <= input(262);
pruneoutput(155) <= input(263);
pruneoutput(156) <= input(264);
pruneoutput(157) <= input(265);
pruneoutput(158) <= input(266);
pruneoutput(159) <= input(267);
pruneoutput(160) <= input(268);
pruneoutput(161) <= input(269);
pruneoutput(162) <= input(270);
pruneoutput(163) <= input(271);
pruneoutput(164) <= input(272);
pruneoutput(165) <= input(273);
pruneoutput(166) <= input(274);
pruneoutput(167) <= input(275);
pruneoutput(168) <= input(276);
pruneoutput(169) <= input(277);
pruneoutput(170) <= input(278);
pruneoutput(171) <= input(279);
pruneoutput(172) <= input(281);
pruneoutput(173) <= input(282);
pruneoutput(174) <= input(283);
pruneoutput(175) <= input(284);
pruneoutput(176) <= input(285);
pruneoutput(177) <= input(286);
pruneoutput(178) <= input(294);
pruneoutput(179) <= input(295);
pruneoutput(180) <= input(296);
pruneoutput(181) <= input(297);
pruneoutput(182) <= input(298);
pruneoutput(183) <= input(299);
pruneoutput(184) <= input(300);
pruneoutput(185) <= input(301);
pruneoutput(186) <= input(302);
pruneoutput(187) <= input(303);
pruneoutput(188) <= input(304);
pruneoutput(189) <= input(305);
pruneoutput(190) <= input(306);
pruneoutput(191) <= input(307);
pruneoutput(192) <= input(309);
pruneoutput(193) <= input(310);
pruneoutput(194) <= input(312);
pruneoutput(195) <= input(313);
pruneoutput(196) <= input(318);
pruneoutput(197) <= input(319);
pruneoutput(198) <= input(320);
pruneoutput(199) <= input(321);
pruneoutput(200) <= input(322);
pruneoutput(201) <= input(323);
pruneoutput(202) <= input(324);
pruneoutput(203) <= input(326);
pruneoutput(204) <= input(327);
pruneoutput(205) <= input(328);
pruneoutput(206) <= input(329);
pruneoutput(207) <= input(330);
pruneoutput(208) <= input(331);
pruneoutput(209) <= input(332);
pruneoutput(210) <= input(333);
pruneoutput(211) <= input(334);
pruneoutput(212) <= input(335);
pruneoutput(213) <= input(336);
pruneoutput(214) <= input(337);
pruneoutput(215) <= input(339);
pruneoutput(216) <= input(340);
pruneoutput(217) <= input(341);
pruneoutput(218) <= input(342);
pruneoutput(219) <= input(346);
pruneoutput(220) <= input(347);
pruneoutput(221) <= input(348);
pruneoutput(222) <= input(349);
pruneoutput(223) <= input(350);
pruneoutput(224) <= input(351);
pruneoutput(225) <= input(352);
pruneoutput(226) <= input(353);
pruneoutput(227) <= input(354);
pruneoutput(228) <= input(355);
pruneoutput(229) <= input(356);
pruneoutput(230) <= input(357);
pruneoutput(231) <= input(358);
pruneoutput(232) <= input(359);
pruneoutput(233) <= input(363);
pruneoutput(234) <= input(364);
pruneoutput(235) <= input(365);
pruneoutput(236) <= input(366);
pruneoutput(237) <= input(367);
pruneoutput(238) <= input(368);
pruneoutput(239) <= input(369);
pruneoutput(240) <= input(370);
pruneoutput(241) <= input(371);
pruneoutput(242) <= input(372);
pruneoutput(243) <= input(373);
pruneoutput(244) <= input(374);
pruneoutput(245) <= input(375);
pruneoutput(246) <= input(376);
pruneoutput(247) <= input(379);
pruneoutput(248) <= input(381);
pruneoutput(249) <= input(382);
pruneoutput(250) <= input(390);
pruneoutput(251) <= input(394);
pruneoutput(252) <= input(395);
pruneoutput(253) <= input(396);
pruneoutput(254) <= input(397);
pruneoutput(255) <= input(398);
pruneoutput(256) <= input(403);
pruneoutput(257) <= input(404);
pruneoutput(258) <= input(405);
pruneoutput(259) <= input(406);
pruneoutput(260) <= input(407);
pruneoutput(261) <= input(408);
pruneoutput(262) <= input(409);
pruneoutput(263) <= input(410);
pruneoutput(264) <= input(411);
pruneoutput(265) <= input(414);
pruneoutput(266) <= input(415);
pruneoutput(267) <= input(418);
pruneoutput(268) <= input(428);
pruneoutput(269) <= input(429);
pruneoutput(270) <= input(430);
pruneoutput(271) <= input(431);
pruneoutput(272) <= input(435);
pruneoutput(273) <= input(441);
pruneoutput(274) <= input(442);
pruneoutput(275) <= input(443);
pruneoutput(276) <= input(447);
pruneoutput(277) <= input(448);
pruneoutput(278) <= input(449);
pruneoutput(279) <= input(450);
pruneoutput(280) <= input(451);
pruneoutput(281) <= input(452);
pruneoutput(282) <= input(454);
pruneoutput(283) <= input(455);
pruneoutput(284) <= input(456);
pruneoutput(285) <= input(457);
pruneoutput(286) <= input(458);
pruneoutput(287) <= input(459);
pruneoutput(288) <= input(465);
pruneoutput(289) <= input(469);
pruneoutput(290) <= input(470);
pruneoutput(291) <= input(471);
pruneoutput(292) <= input(472);
pruneoutput(293) <= input(473);
pruneoutput(294) <= input(478);
pruneoutput(295) <= input(479);
pruneoutput(296) <= input(480);
pruneoutput(297) <= input(482);
pruneoutput(298) <= input(487);
pruneoutput(299) <= input(488);
pruneoutput(300) <= input(489);
pruneoutput(301) <= input(490);
pruneoutput(302) <= input(491);
pruneoutput(303) <= input(492);
pruneoutput(304) <= input(493);
pruneoutput(305) <= input(494);
pruneoutput(306) <= input(495);
pruneoutput(307) <= input(496);
pruneoutput(308) <= input(497);
pruneoutput(309) <= input(498);
pruneoutput(310) <= input(500);
pruneoutput(311) <= input(501);
pruneoutput(312) <= input(502);
pruneoutput(313) <= input(503);
pruneoutput(314) <= input(504);
pruneoutput(315) <= input(505);
pruneoutput(316) <= input(506);
pruneoutput(317) <= input(507);
pruneoutput(318) <= input(508);
pruneoutput(319) <= input(509);
pruneoutput(320) <= input(510);
pruneoutput(321) <= input(511);
pruneoutput(322) <= input(512);
pruneoutput(323) <= input(513);
pruneoutput(324) <= input(514);
pruneoutput(325) <= input(515);
pruneoutput(326) <= input(516);
pruneoutput(327) <= input(517);
pruneoutput(328) <= input(518);
pruneoutput(329) <= input(519);
pruneoutput(330) <= input(520);
pruneoutput(331) <= input(521);
pruneoutput(332) <= input(522);
pruneoutput(333) <= input(523);
pruneoutput(334) <= input(524);
pruneoutput(335) <= input(525);
pruneoutput(336) <= input(526);
pruneoutput(337) <= input(527);
pruneoutput(338) <= input(528);
pruneoutput(339) <= input(530);
pruneoutput(340) <= input(531);
pruneoutput(341) <= input(537);
pruneoutput(342) <= input(538);
pruneoutput(343) <= input(539);
pruneoutput(344) <= input(540);
pruneoutput(345) <= input(541);
pruneoutput(346) <= input(542);
pruneoutput(347) <= input(543);
pruneoutput(348) <= input(544);
pruneoutput(349) <= input(545);
pruneoutput(350) <= input(547);
pruneoutput(351) <= input(551);
pruneoutput(352) <= input(552);
pruneoutput(353) <= input(553);
pruneoutput(354) <= input(554);
pruneoutput(355) <= input(555);
pruneoutput(356) <= input(556);
pruneoutput(357) <= input(557);
pruneoutput(358) <= input(558);
pruneoutput(359) <= input(559);
pruneoutput(360) <= input(560);
pruneoutput(361) <= input(561);
pruneoutput(362) <= input(562);
pruneoutput(363) <= input(563);
pruneoutput(364) <= input(565);
pruneoutput(365) <= input(566);
pruneoutput(366) <= input(567);
pruneoutput(367) <= input(568);
pruneoutput(368) <= input(569);
pruneoutput(369) <= input(570);
pruneoutput(370) <= input(571);
pruneoutput(371) <= input(572);
pruneoutput(372) <= input(573);
pruneoutput(373) <= input(574);
pruneoutput(374) <= input(575);
pruneoutput(375) <= input(576);
pruneoutput(376) <= input(577);
pruneoutput(377) <= input(578);
pruneoutput(378) <= input(579);
pruneoutput(379) <= input(583);
pruneoutput(380) <= input(586);
pruneoutput(381) <= input(588);
pruneoutput(382) <= input(589);
pruneoutput(383) <= input(596);
pruneoutput(384) <= input(597);
pruneoutput(385) <= input(598);
pruneoutput(386) <= input(599);
pruneoutput(387) <= input(600);
pruneoutput(388) <= input(601);
pruneoutput(389) <= input(603);
pruneoutput(390) <= input(604);
pruneoutput(391) <= input(605);
pruneoutput(392) <= input(606);
pruneoutput(393) <= input(607);
pruneoutput(394) <= input(608);
pruneoutput(395) <= input(609);
pruneoutput(396) <= input(610);
pruneoutput(397) <= input(611);
pruneoutput(398) <= input(612);
pruneoutput(399) <= input(613);
pruneoutput(400) <= input(614);
pruneoutput(401) <= input(615);
pruneoutput(402) <= input(616);
pruneoutput(403) <= input(617);
pruneoutput(404) <= input(618);
pruneoutput(405) <= input(623);
pruneoutput(406) <= input(625);
pruneoutput(407) <= input(626);
pruneoutput(408) <= input(627);
pruneoutput(409) <= input(628);
pruneoutput(410) <= input(637);
pruneoutput(411) <= input(638);
pruneoutput(412) <= input(639);
pruneoutput(413) <= input(642);
pruneoutput(414) <= input(644);
pruneoutput(415) <= input(645);
pruneoutput(416) <= input(646);
pruneoutput(417) <= input(647);
pruneoutput(418) <= input(648);
pruneoutput(419) <= input(649);
pruneoutput(420) <= input(650);
pruneoutput(421) <= input(651);
pruneoutput(422) <= input(652);
pruneoutput(423) <= input(659);
pruneoutput(424) <= input(660);
pruneoutput(425) <= input(661);
pruneoutput(426) <= input(662);
pruneoutput(427) <= input(663);
pruneoutput(428) <= input(664);
pruneoutput(429) <= input(665);
pruneoutput(430) <= input(666);
pruneoutput(431) <= input(667);
pruneoutput(432) <= input(668);
pruneoutput(433) <= input(669);
pruneoutput(434) <= input(670);
pruneoutput(435) <= input(671);
pruneoutput(436) <= input(672);
pruneoutput(437) <= input(673);
pruneoutput(438) <= input(674);
pruneoutput(439) <= input(675);
pruneoutput(440) <= input(676);
pruneoutput(441) <= input(677);
pruneoutput(442) <= input(678);
pruneoutput(443) <= input(679);
pruneoutput(444) <= input(680);
pruneoutput(445) <= input(684);
pruneoutput(446) <= input(685);
pruneoutput(447) <= input(686);
pruneoutput(448) <= input(687);
pruneoutput(449) <= input(689);
pruneoutput(450) <= input(690);
pruneoutput(451) <= input(691);
pruneoutput(452) <= input(692);
pruneoutput(453) <= input(695);
pruneoutput(454) <= input(696);
pruneoutput(455) <= input(697);
pruneoutput(456) <= input(698);
pruneoutput(457) <= input(699);
pruneoutput(458) <= input(702);
pruneoutput(459) <= input(703);
pruneoutput(460) <= input(704);
pruneoutput(461) <= input(705);
pruneoutput(462) <= input(706);
pruneoutput(463) <= input(707);
pruneoutput(464) <= input(709);
pruneoutput(465) <= input(710);
pruneoutput(466) <= input(712);
pruneoutput(467) <= input(713);
pruneoutput(468) <= input(714);
pruneoutput(469) <= input(722);
pruneoutput(470) <= input(723);
pruneoutput(471) <= input(724);
pruneoutput(472) <= input(725);
pruneoutput(473) <= input(726);
pruneoutput(474) <= input(727);
pruneoutput(475) <= input(728);
pruneoutput(476) <= input(730);
pruneoutput(477) <= input(731);
pruneoutput(478) <= input(732);
pruneoutput(479) <= input(737);
pruneoutput(480) <= input(738);
pruneoutput(481) <= input(739);
pruneoutput(482) <= input(743);
pruneoutput(483) <= input(744);
pruneoutput(484) <= input(745);
pruneoutput(485) <= input(746);
pruneoutput(486) <= input(747);
pruneoutput(487) <= input(748);
pruneoutput(488) <= input(749);
pruneoutput(489) <= input(750);
pruneoutput(490) <= input(751);
pruneoutput(491) <= input(752);
pruneoutput(492) <= input(753);
pruneoutput(493) <= input(754);
pruneoutput(494) <= input(755);
pruneoutput(495) <= input(756);
pruneoutput(496) <= input(757);
pruneoutput(497) <= input(758);
pruneoutput(498) <= input(759);
pruneoutput(499) <= input(760);
pruneoutput(500) <= input(761);
pruneoutput(501) <= input(765);
pruneoutput(502) <= input(767);
pruneoutput(503) <= input(768);
pruneoutput(504) <= input(769);
pruneoutput(505) <= input(770);
pruneoutput(506) <= input(771);
pruneoutput(507) <= input(772);
pruneoutput(508) <= input(774);
pruneoutput(509) <= input(775);
pruneoutput(510) <= input(776);
pruneoutput(511) <= input(778);
pruneoutput(512) <= input(779);
pruneoutput(513) <= input(781);
pruneoutput(514) <= input(782);
pruneoutput(515) <= input(783);
pruneoutput(516) <= input(784);
pruneoutput(517) <= input(785);
pruneoutput(518) <= input(786);
pruneoutput(519) <= input(787);
pruneoutput(520) <= input(788);
pruneoutput(521) <= input(789);
pruneoutput(522) <= input(790);
pruneoutput(523) <= input(791);
pruneoutput(524) <= input(792);
pruneoutput(525) <= input(793);
pruneoutput(526) <= input(794);
pruneoutput(527) <= input(795);
pruneoutput(528) <= input(796);
pruneoutput(529) <= input(797);
pruneoutput(530) <= input(798);
pruneoutput(531) <= input(799);
pruneoutput(532) <= input(804);
pruneoutput(533) <= input(805);
pruneoutput(534) <= input(806);
pruneoutput(535) <= input(807);
pruneoutput(536) <= input(808);
pruneoutput(537) <= input(809);
pruneoutput(538) <= input(810);
pruneoutput(539) <= input(811);
pruneoutput(540) <= input(813);
pruneoutput(541) <= input(814);
pruneoutput(542) <= input(815);
pruneoutput(543) <= input(816);
pruneoutput(544) <= input(817);
pruneoutput(545) <= input(818);
pruneoutput(546) <= input(822);
pruneoutput(547) <= input(823);
pruneoutput(548) <= input(824);
pruneoutput(549) <= input(825);
pruneoutput(550) <= input(829);
pruneoutput(551) <= input(830);
pruneoutput(552) <= input(831);
pruneoutput(553) <= input(832);
pruneoutput(554) <= input(833);
pruneoutput(555) <= input(834);
pruneoutput(556) <= input(835);
pruneoutput(557) <= input(836);
pruneoutput(558) <= input(843);
pruneoutput(559) <= input(852);
pruneoutput(560) <= input(853);
pruneoutput(561) <= input(854);
pruneoutput(562) <= input(856);
pruneoutput(563) <= input(857);
pruneoutput(564) <= input(858);
pruneoutput(565) <= input(859);
pruneoutput(566) <= input(860);
pruneoutput(567) <= input(861);
pruneoutput(568) <= input(864);
pruneoutput(569) <= input(869);
pruneoutput(570) <= input(870);
pruneoutput(571) <= input(878);
pruneoutput(572) <= input(879);
pruneoutput(573) <= input(882);
pruneoutput(574) <= input(883);
pruneoutput(575) <= input(884);
pruneoutput(576) <= input(885);
pruneoutput(577) <= input(886);
pruneoutput(578) <= input(887);
pruneoutput(579) <= input(888);
pruneoutput(580) <= input(892);
pruneoutput(581) <= input(894);
pruneoutput(582) <= input(895);
pruneoutput(583) <= input(896);
pruneoutput(584) <= input(897);
pruneoutput(585) <= input(898);
pruneoutput(586) <= input(899);
pruneoutput(587) <= input(902);
pruneoutput(588) <= input(903);
pruneoutput(589) <= input(904);
pruneoutput(590) <= input(905);
pruneoutput(591) <= input(906);
pruneoutput(592) <= input(907);
pruneoutput(593) <= input(908);
pruneoutput(594) <= input(909);
pruneoutput(595) <= input(915);
pruneoutput(596) <= input(916);
pruneoutput(597) <= input(917);
pruneoutput(598) <= input(929);
pruneoutput(599) <= input(930);
pruneoutput(600) <= input(931);
pruneoutput(601) <= input(934);
pruneoutput(602) <= input(935);
pruneoutput(603) <= input(936);
pruneoutput(604) <= input(938);
pruneoutput(605) <= input(939);
pruneoutput(606) <= input(940);
pruneoutput(607) <= input(941);
pruneoutput(608) <= input(942);
pruneoutput(609) <= input(943);
pruneoutput(610) <= input(944);
pruneoutput(611) <= input(945);
pruneoutput(612) <= input(946);
pruneoutput(613) <= input(947);
pruneoutput(614) <= input(948);
pruneoutput(615) <= input(949);
pruneoutput(616) <= input(950);
pruneoutput(617) <= input(951);
pruneoutput(618) <= input(952);
pruneoutput(619) <= input(953);
pruneoutput(620) <= input(954);
pruneoutput(621) <= input(956);
pruneoutput(622) <= input(957);
pruneoutput(623) <= input(958);
pruneoutput(624) <= input(962);
pruneoutput(625) <= input(963);
pruneoutput(626) <= input(964);
pruneoutput(627) <= input(966);
pruneoutput(628) <= input(968);
pruneoutput(629) <= input(971);
pruneoutput(630) <= input(973);
pruneoutput(631) <= input(974);
pruneoutput(632) <= input(975);
pruneoutput(633) <= input(976);
pruneoutput(634) <= input(979);
pruneoutput(635) <= input(980);
pruneoutput(636) <= input(981);
pruneoutput(637) <= input(982);
pruneoutput(638) <= input(983);
pruneoutput(639) <= input(984);
pruneoutput(640) <= input(988);
pruneoutput(641) <= input(989);
pruneoutput(642) <= input(990);
pruneoutput(643) <= input(991);
pruneoutput(644) <= input(992);
pruneoutput(645) <= input(994);

END ARCHITECTURE behavioral;