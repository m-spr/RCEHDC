-- MIT License

-- Copyright (c) 2024 m-spr

-- Permission is hereby granted, free of charge, to any person obtaining a copy
-- of this software and associated documentation files (the "Software"), to deal
-- in the Software without restriction, including without limitation the rights
-- to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
-- copies of the Software, and to permit persons to whom the Software is
-- furnished to do so, subject to the following conditions:

-- The above copyright notice and this permission notice shall be included in all
-- copies or substantial portions of the Software.

-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
-- IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
-- FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
-- AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
-- LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
-- OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
-- SOFTWARE.

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY BasedVectorLFSR IS
    GENERIC (
        n : INTEGER := 2000  -- Number of bits
    );	 
    PORT (
        clk  : IN STD_LOGIC;
        rst  : IN STD_LOGIC;
        update : IN STD_LOGIC; 
        congigSignitureIn  : IN STD_LOGIC_VECTOR (n-1 DOWNTO 0);
        congigInitialvaluesIn : IN STD_LOGIC_VECTOR (n-1 DOWNTO 0);
        dout : OUT STD_LOGIC_VECTOR (n-1 DOWNTO 0)
    );
END ENTITY BasedVectorLFSR;

ARCHITECTURE behavioral OF BasedVectorLFSR IS

    COMPONENT regOne IS
        GENERIC (
            init : STD_LOGIC := '1'  -- Initial value
        );
        PORT (
            clk       : IN STD_LOGIC;
            regUpdate : IN STD_LOGIC;
            regrst    : IN STD_LOGIC;
            din       : IN STD_LOGIC;
            dout      : OUT STD_LOGIC
        );
    END COMPONENT;

    SIGNAL interValIn, interValOut : STD_LOGIC_VECTOR (n-1 DOWNTO 0);
    SIGNAL interValOutR : STD_LOGIC_VECTOR (0 TO n-1);

    CONSTANT congigSigniture : STD_LOGIC_VECTOR (n-1 DOWNTO 0) :=    "1100011001101000001010100111100110101010000110110101010000010010111010000000001001101011000011111100100010011111111110101100010101110101000011101111111101101100111011000001001011111011100000110101001011101000101001011110011000111101001100100100011100101001000000001011010101000110001100101001001011101101110110111010101010101001100001110011010001001110010010010111010000000010010111011110101010010111101101010110100000001101101011011011000001011000010111110111010010111000000011110001010001110101110010001011010010000010000010000010001001001001110101100111011010010110000011011000101010100110000101101011011101111000011001000110101110101011010010111000101010010000100101100100101000010000110100000100111001110111110001111100001110101011100001100111101000000110100010011110001001111000010001001011100010111010110010001000001000001001111000111001010110011111001010100101001101011000111001010010011100100101011100111000001100100101000111011110110100010011011000100111000000110000101011110111010000001011"; 

    CONSTANT congigInitialvalues : STD_LOGIC_VECTOR (n-1 DOWNTO 0) := "1100011111100001110000010001110000100000101101000111010010010010110001011101100001100010001111100001111110000011110110000111100001011110111110010011110011100101101010100110001010100101110100111001101100011100110111010000010111011111011101001001111001111110001000010011000000111101100111101001111101111010101010001001000111111110101001011000101010010101011010110100000011110110000111100100110101101111101100110010011010001101010100011011001000011000100100010110110000000010000001000100101111111000101001101000000101111010100100011110001011001101110000011011001110011010110101101111010100010011100010010000000101010001011100101000101010010000110110000000000110010110100011000010111010010011011001101001100000100101001000100000100010000000111011110110111101000110001101001010110100011100111111001110110001100000101000100111101001111101011000100000010100100001110000110100011111011100010010101001100101010110101011011011000010010001101100001011011100110100011110110000001001100011111100111100110111111010";

BEGIN

    -- Generate Registers
    regArr : FOR i IN 1 TO n-1 GENERATE
        Ireg : regOne 
            GENERIC MAP (congigInitialvalues(i))
            PORT MAP (
                clk      => clk,  
                regUpdate => update, 
                regrst   => rst, 
                din      => interValIn(i),  
                dout     => interValOut(i) 
            );   
    END GENERATE regArr;

    -- Generate XOR Chain
    xorchain : FOR i IN 1 TO n-1 GENERATE
        xorchain1: IF (congigSigniture(i) = '1') GENERATE
            interValIn(i) <= interValOut(i-1) XOR interValOut(n-1);
        END GENERATE xorchain1;

        xorchain2: IF (congigSigniture(i) = '0') GENERATE
            interValIn(i) <= interValOut(i-1);
        END GENERATE xorchain2;
    END GENERATE xorchain;

    -- First Register
    interValIn(0) <= interValOut(n-1);
    
    reg0 : regOne 
        GENERIC MAP (congigInitialvalues(0))
        PORT MAP (
            clk      => clk,  
            regUpdate => update, 
            regrst   => rst, 
            din      => interValIn(0),  
            dout     => interValOut(0)
        ); 

    -- Output Assignment
    dout <= interValOut;

END ARCHITECTURE behavioral;
