LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY BasedVectorLFSR IS
	GENERIC ( n	: INTEGER	:= 2000			    -- number of bits
				);	 
	PORT (
		clk, rst, update	: IN STD_LOGIC; 
		congigSignitureIn , congigInitialvaluesIn : IN STD_LOGIC_VECTOR (n-1 DOWNTO 0 );
		dout				: OUT  STD_LOGIC_VECTOR (n-1 DOWNTO 0 )
	);
END ENTITY BasedVectorLFSR;

ARCHITECTURE behavioral OF BasedVectorLFSR IS

COMPONENT  regOne IS
	GENERIC (init : STD_LOGIC := '1');   -- initial value
	PORT (
		clk 				: IN  STD_LOGIC;
		regUpdate, regrst 	: IN  STD_LOGIC;
		din        			: IN  STD_LOGIC;
		dout        		: OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL interValIn : STD_LOGIC_VECTOR (n-1 DOWNTO 0);
SIGNAL interValOut : STD_LOGIC_VECTOR (n-1 DOWNTO 0);
SIGNAL interValOutR : STD_LOGIC_VECTOR (0 TO n-1);
CONSTANT congigSigniture : STD_LOGIC_VECTOR (n-1 DOWNTO 0) :=    "1101101001001100101111100000110011000000011111011101000011110011010101110001001011100000010000000100011100011011111100110100010010001001100010011101101011010110101001000000010010010011011111110001100011010011110011011110111001100000111110101101000001100001010011110011111010100000001100110010110001010100101100111001101000010001001000011010110111010011001111101101100110010011110011000001001101001010110000101011111101010000011100001010100101001010110001011101101000101010110010000010001001010110100101000101010111000010000100000011110000110110111111110001100100001011011111111101100111001111001011100100000000010111010111101110000011000000111100100101111001101001100001101000000000111001010111010001000001101101101010101101000011110010011000111110110110000010111011010110001111101110001101100110011010100011001110001010001010000000000010101000101010011000110100110100001101110111011111001101111110111110101010111011001010001011111101000100000101000011111010110001010001000111110100011100011100000000"; --"1010101011000011001011001000001001000110100100000010011011000001110101100010000001000111100011101100011001100110100010101100010001011111010110000011000010111011110110101000110101100100110110100001010010111100101010101000111011111101101111011111001111001010110000010110100001111110011100100000000110110110000000011011010111101011100110101100010100100011010011000001010111000000010001101101101011010110110011110000010000110110010110100011111001011110011010011101011010111100011001010111011111110101100110001110000011111111110110001011001111111110010101010010011101000011100111101011011000110101010101100000100001101010101000111111001001111101010000110001110110001010111000101100101010011110010101100010011011011111111100100111100010011100101010010000001100111011100101101011100010111001000110101111110111111010001000100101100011100010001011001100110111011010101010000010100000000101001000110011011011011100010011011001001011100000000000000001000010010101100101110110001001101010101101010001110000001100";

CONSTANT congigInitialvalues : STD_LOGIC_VECTOR (n-1 DOWNTO 0) := "1001100110010010100011010110111010001010010100001000100000000110101011001110100001011101000101000100001001011001111111101111100101100000001010111001111110101110101011111001010101110110111000100110110101110101010111011000010010101011101101100101001010110010000010100110100000100111011110010100111101100111000000011000010011000110100000010000110110111011010001101001100100110000110010010010000110001111000101010100010001011101011001010111100100100110111001110110001001011101101011000001010110111101111100111011011001001100010000110000011111100110101001010110111100000101000010011101101010111001100001111011001011100001111011010000011000110111100000111110001001101110110011000010111101110110010000000011110111100011111000000100011100000011000110001110101110101100000111000100100110101111100100101011111111000010011000100101111100100110110001001110011010100100001101010010100110100110001101000100101111110110101000011011010101010000110100001001001001110000100010001101001010101100101000010011001100010010";--"1111000000100110110100000110111010000101111100010011000110000110000100100100100010111110100100111000000001010111001001001000111010011010000001011010010100111000100010110111010111110010000101010100011101011111011100001011010100011100110110100001101100111100101111001001100100000011110111000110111000010001111100011110001110001010001011011011000000001010000001000001000011100010110011111101111000000010000111110001101011110111101010101010001110110110100100101011011011011110000111110110011000100110111010000011101100111010000010101011010111001011110110100000101100101111110011010011010010111000100100101100101101010001001110100010100001011100010111110010110011101000111110110001100100011100001110110000101111110011100100011011011101101110010101000101010100101011110011100100111100010011011100100101001010000110000101011100001110011111100011000011101010100001011010100101011110000100010001101001000000001011010001001001001000111010110101000010101011111110000010001010100111111100100011000110110101100110";

BEGIN

	regArr : FOR i IN 1 TO n-1 GENERATE
		Ireg : regOne 
			GENERIC map(congigInitialvalues(i))
			PORT map(clk,  update, rst, 
			interValIn(i), 	interValOut(i) 
					 );   
	END GENERATE regArr;
	xorchain : FOR i IN 1 TO n-1 GENERATE
	xorchain1: IF (congigSigniture(i) = '1') GENERATE
			interValIn(i) <= interValOut(i-1) XOR  interValOut(n-1);
		END GENERATE xorchain1;
	xorchain2: IF (congigSigniture(i) = '0') GENERATE
			interValIn(i) <= interValOut(i-1);
		END GENERATE xorchain2;
	END GENERATE xorchain;
	interValIn(0) <= interValOut(n-1);
	reg0 : regOne 
			GENERIC map(congigInitialvalues(0))
			PORT map(clk,  update, rst, 
			interValIn(0), 	interValOut(0) 
					 ); 
	--interValOutR <= interValOut;
	dout <= interValOut;--(0 TO n-1);

END ARCHITECTURE behavioral;