LIBRARY IEEE; 
USE IEEE.STD_LOGIC_1164.ALL; 
USE IEEE.NUMERIC_STD.ALL; 
  
ENTITY connector IS 
	PORT ( 
		input         : IN  STD_LOGIC_VECTOR (999 DOWNTO 0); 
		pruneoutput        : OUT  STD_LOGIC_VECTOR (640 DOWNTO 0)      
	);
END ENTITY connector;

ARCHITECTURE behavioral OF connector  IS
BEGIN
pruneoutput(0) <= input(0);
pruneoutput(1) <= input(1);
pruneoutput(2) <= input(2);
pruneoutput(3) <= input(3);
pruneoutput(4) <= input(4);
pruneoutput(5) <= input(7);
pruneoutput(6) <= input(8);
pruneoutput(7) <= input(9);
pruneoutput(8) <= input(11);
pruneoutput(9) <= input(14);
pruneoutput(10) <= input(15);
pruneoutput(11) <= input(16);
pruneoutput(12) <= input(17);
pruneoutput(13) <= input(18);
pruneoutput(14) <= input(19);
pruneoutput(15) <= input(20);
pruneoutput(16) <= input(21);
pruneoutput(17) <= input(22);
pruneoutput(18) <= input(23);
pruneoutput(19) <= input(24);
pruneoutput(20) <= input(25);
pruneoutput(21) <= input(26);
pruneoutput(22) <= input(27);
pruneoutput(23) <= input(28);
pruneoutput(24) <= input(29);
pruneoutput(25) <= input(30);
pruneoutput(26) <= input(34);
pruneoutput(27) <= input(35);
pruneoutput(28) <= input(36);
pruneoutput(29) <= input(37);
pruneoutput(30) <= input(38);
pruneoutput(31) <= input(40);
pruneoutput(32) <= input(41);
pruneoutput(33) <= input(42);
pruneoutput(34) <= input(43);
pruneoutput(35) <= input(51);
pruneoutput(36) <= input(52);
pruneoutput(37) <= input(53);
pruneoutput(38) <= input(54);
pruneoutput(39) <= input(55);
pruneoutput(40) <= input(56);
pruneoutput(41) <= input(58);
pruneoutput(42) <= input(59);
pruneoutput(43) <= input(60);
pruneoutput(44) <= input(61);
pruneoutput(45) <= input(62);
pruneoutput(46) <= input(63);
pruneoutput(47) <= input(66);
pruneoutput(48) <= input(67);
pruneoutput(49) <= input(75);
pruneoutput(50) <= input(76);
pruneoutput(51) <= input(77);
pruneoutput(52) <= input(78);
pruneoutput(53) <= input(79);
pruneoutput(54) <= input(80);
pruneoutput(55) <= input(81);
pruneoutput(56) <= input(84);
pruneoutput(57) <= input(85);
pruneoutput(58) <= input(86);
pruneoutput(59) <= input(87);
pruneoutput(60) <= input(89);
pruneoutput(61) <= input(90);
pruneoutput(62) <= input(91);
pruneoutput(63) <= input(92);
pruneoutput(64) <= input(94);
pruneoutput(65) <= input(97);
pruneoutput(66) <= input(101);
pruneoutput(67) <= input(102);
pruneoutput(68) <= input(107);
pruneoutput(69) <= input(108);
pruneoutput(70) <= input(109);
pruneoutput(71) <= input(111);
pruneoutput(72) <= input(112);
pruneoutput(73) <= input(113);
pruneoutput(74) <= input(114);
pruneoutput(75) <= input(115);
pruneoutput(76) <= input(116);
pruneoutput(77) <= input(117);
pruneoutput(78) <= input(118);
pruneoutput(79) <= input(121);
pruneoutput(80) <= input(122);
pruneoutput(81) <= input(123);
pruneoutput(82) <= input(124);
pruneoutput(83) <= input(125);
pruneoutput(84) <= input(126);
pruneoutput(85) <= input(127);
pruneoutput(86) <= input(128);
pruneoutput(87) <= input(129);
pruneoutput(88) <= input(132);
pruneoutput(89) <= input(133);
pruneoutput(90) <= input(134);
pruneoutput(91) <= input(135);
pruneoutput(92) <= input(136);
pruneoutput(93) <= input(137);
pruneoutput(94) <= input(148);
pruneoutput(95) <= input(149);
pruneoutput(96) <= input(150);
pruneoutput(97) <= input(151);
pruneoutput(98) <= input(152);
pruneoutput(99) <= input(153);
pruneoutput(100) <= input(154);
pruneoutput(101) <= input(156);
pruneoutput(102) <= input(159);
pruneoutput(103) <= input(162);
pruneoutput(104) <= input(163);
pruneoutput(105) <= input(164);
pruneoutput(106) <= input(165);
pruneoutput(107) <= input(166);
pruneoutput(108) <= input(167);
pruneoutput(109) <= input(168);
pruneoutput(110) <= input(171);
pruneoutput(111) <= input(172);
pruneoutput(112) <= input(173);
pruneoutput(113) <= input(174);
pruneoutput(114) <= input(175);
pruneoutput(115) <= input(179);
pruneoutput(116) <= input(180);
pruneoutput(117) <= input(181);
pruneoutput(118) <= input(185);
pruneoutput(119) <= input(186);
pruneoutput(120) <= input(187);
pruneoutput(121) <= input(188);
pruneoutput(122) <= input(189);
pruneoutput(123) <= input(190);
pruneoutput(124) <= input(196);
pruneoutput(125) <= input(197);
pruneoutput(126) <= input(201);
pruneoutput(127) <= input(202);
pruneoutput(128) <= input(203);
pruneoutput(129) <= input(206);
pruneoutput(130) <= input(207);
pruneoutput(131) <= input(208);
pruneoutput(132) <= input(211);
pruneoutput(133) <= input(212);
pruneoutput(134) <= input(215);
pruneoutput(135) <= input(221);
pruneoutput(136) <= input(222);
pruneoutput(137) <= input(223);
pruneoutput(138) <= input(224);
pruneoutput(139) <= input(225);
pruneoutput(140) <= input(232);
pruneoutput(141) <= input(233);
pruneoutput(142) <= input(234);
pruneoutput(143) <= input(235);
pruneoutput(144) <= input(236);
pruneoutput(145) <= input(238);
pruneoutput(146) <= input(239);
pruneoutput(147) <= input(240);
pruneoutput(148) <= input(242);
pruneoutput(149) <= input(243);
pruneoutput(150) <= input(244);
pruneoutput(151) <= input(245);
pruneoutput(152) <= input(246);
pruneoutput(153) <= input(247);
pruneoutput(154) <= input(249);
pruneoutput(155) <= input(250);
pruneoutput(156) <= input(251);
pruneoutput(157) <= input(252);
pruneoutput(158) <= input(253);
pruneoutput(159) <= input(254);
pruneoutput(160) <= input(255);
pruneoutput(161) <= input(256);
pruneoutput(162) <= input(257);
pruneoutput(163) <= input(258);
pruneoutput(164) <= input(259);
pruneoutput(165) <= input(260);
pruneoutput(166) <= input(261);
pruneoutput(167) <= input(262);
pruneoutput(168) <= input(263);
pruneoutput(169) <= input(264);
pruneoutput(170) <= input(265);
pruneoutput(171) <= input(266);
pruneoutput(172) <= input(267);
pruneoutput(173) <= input(268);
pruneoutput(174) <= input(269);
pruneoutput(175) <= input(270);
pruneoutput(176) <= input(271);
pruneoutput(177) <= input(272);
pruneoutput(178) <= input(273);
pruneoutput(179) <= input(275);
pruneoutput(180) <= input(276);
pruneoutput(181) <= input(277);
pruneoutput(182) <= input(278);
pruneoutput(183) <= input(280);
pruneoutput(184) <= input(281);
pruneoutput(185) <= input(283);
pruneoutput(186) <= input(286);
pruneoutput(187) <= input(287);
pruneoutput(188) <= input(288);
pruneoutput(189) <= input(292);
pruneoutput(190) <= input(293);
pruneoutput(191) <= input(294);
pruneoutput(192) <= input(295);
pruneoutput(193) <= input(299);
pruneoutput(194) <= input(303);
pruneoutput(195) <= input(311);
pruneoutput(196) <= input(313);
pruneoutput(197) <= input(314);
pruneoutput(198) <= input(315);
pruneoutput(199) <= input(316);
pruneoutput(200) <= input(317);
pruneoutput(201) <= input(318);
pruneoutput(202) <= input(319);
pruneoutput(203) <= input(320);
pruneoutput(204) <= input(321);
pruneoutput(205) <= input(323);
pruneoutput(206) <= input(324);
pruneoutput(207) <= input(325);
pruneoutput(208) <= input(326);
pruneoutput(209) <= input(330);
pruneoutput(210) <= input(331);
pruneoutput(211) <= input(332);
pruneoutput(212) <= input(337);
pruneoutput(213) <= input(338);
pruneoutput(214) <= input(339);
pruneoutput(215) <= input(340);
pruneoutput(216) <= input(341);
pruneoutput(217) <= input(347);
pruneoutput(218) <= input(348);
pruneoutput(219) <= input(349);
pruneoutput(220) <= input(350);
pruneoutput(221) <= input(351);
pruneoutput(222) <= input(352);
pruneoutput(223) <= input(353);
pruneoutput(224) <= input(354);
pruneoutput(225) <= input(355);
pruneoutput(226) <= input(356);
pruneoutput(227) <= input(357);
pruneoutput(228) <= input(363);
pruneoutput(229) <= input(365);
pruneoutput(230) <= input(366);
pruneoutput(231) <= input(367);
pruneoutput(232) <= input(370);
pruneoutput(233) <= input(373);
pruneoutput(234) <= input(374);
pruneoutput(235) <= input(375);
pruneoutput(236) <= input(376);
pruneoutput(237) <= input(377);
pruneoutput(238) <= input(378);
pruneoutput(239) <= input(379);
pruneoutput(240) <= input(380);
pruneoutput(241) <= input(381);
pruneoutput(242) <= input(382);
pruneoutput(243) <= input(383);
pruneoutput(244) <= input(384);
pruneoutput(245) <= input(386);
pruneoutput(246) <= input(387);
pruneoutput(247) <= input(388);
pruneoutput(248) <= input(391);
pruneoutput(249) <= input(392);
pruneoutput(250) <= input(393);
pruneoutput(251) <= input(394);
pruneoutput(252) <= input(395);
pruneoutput(253) <= input(399);
pruneoutput(254) <= input(400);
pruneoutput(255) <= input(401);
pruneoutput(256) <= input(406);
pruneoutput(257) <= input(413);
pruneoutput(258) <= input(414);
pruneoutput(259) <= input(418);
pruneoutput(260) <= input(419);
pruneoutput(261) <= input(420);
pruneoutput(262) <= input(421);
pruneoutput(263) <= input(424);
pruneoutput(264) <= input(425);
pruneoutput(265) <= input(435);
pruneoutput(266) <= input(436);
pruneoutput(267) <= input(437);
pruneoutput(268) <= input(438);
pruneoutput(269) <= input(439);
pruneoutput(270) <= input(440);
pruneoutput(271) <= input(441);
pruneoutput(272) <= input(442);
pruneoutput(273) <= input(443);
pruneoutput(274) <= input(444);
pruneoutput(275) <= input(445);
pruneoutput(276) <= input(446);
pruneoutput(277) <= input(447);
pruneoutput(278) <= input(448);
pruneoutput(279) <= input(449);
pruneoutput(280) <= input(450);
pruneoutput(281) <= input(453);
pruneoutput(282) <= input(454);
pruneoutput(283) <= input(455);
pruneoutput(284) <= input(457);
pruneoutput(285) <= input(458);
pruneoutput(286) <= input(459);
pruneoutput(287) <= input(460);
pruneoutput(288) <= input(461);
pruneoutput(289) <= input(462);
pruneoutput(290) <= input(465);
pruneoutput(291) <= input(466);
pruneoutput(292) <= input(471);
pruneoutput(293) <= input(472);
pruneoutput(294) <= input(473);
pruneoutput(295) <= input(475);
pruneoutput(296) <= input(476);
pruneoutput(297) <= input(477);
pruneoutput(298) <= input(478);
pruneoutput(299) <= input(479);
pruneoutput(300) <= input(480);
pruneoutput(301) <= input(481);
pruneoutput(302) <= input(482);
pruneoutput(303) <= input(484);
pruneoutput(304) <= input(485);
pruneoutput(305) <= input(486);
pruneoutput(306) <= input(487);
pruneoutput(307) <= input(488);
pruneoutput(308) <= input(489);
pruneoutput(309) <= input(490);
pruneoutput(310) <= input(493);
pruneoutput(311) <= input(496);
pruneoutput(312) <= input(497);
pruneoutput(313) <= input(500);
pruneoutput(314) <= input(501);
pruneoutput(315) <= input(502);
pruneoutput(316) <= input(503);
pruneoutput(317) <= input(504);
pruneoutput(318) <= input(506);
pruneoutput(319) <= input(511);
pruneoutput(320) <= input(512);
pruneoutput(321) <= input(515);
pruneoutput(322) <= input(516);
pruneoutput(323) <= input(519);
pruneoutput(324) <= input(520);
pruneoutput(325) <= input(522);
pruneoutput(326) <= input(523);
pruneoutput(327) <= input(525);
pruneoutput(328) <= input(526);
pruneoutput(329) <= input(527);
pruneoutput(330) <= input(528);
pruneoutput(331) <= input(529);
pruneoutput(332) <= input(530);
pruneoutput(333) <= input(531);
pruneoutput(334) <= input(538);
pruneoutput(335) <= input(541);
pruneoutput(336) <= input(543);
pruneoutput(337) <= input(544);
pruneoutput(338) <= input(545);
pruneoutput(339) <= input(548);
pruneoutput(340) <= input(549);
pruneoutput(341) <= input(553);
pruneoutput(342) <= input(554);
pruneoutput(343) <= input(555);
pruneoutput(344) <= input(556);
pruneoutput(345) <= input(557);
pruneoutput(346) <= input(558);
pruneoutput(347) <= input(559);
pruneoutput(348) <= input(560);
pruneoutput(349) <= input(561);
pruneoutput(350) <= input(562);
pruneoutput(351) <= input(563);
pruneoutput(352) <= input(564);
pruneoutput(353) <= input(565);
pruneoutput(354) <= input(566);
pruneoutput(355) <= input(567);
pruneoutput(356) <= input(569);
pruneoutput(357) <= input(570);
pruneoutput(358) <= input(571);
pruneoutput(359) <= input(572);
pruneoutput(360) <= input(573);
pruneoutput(361) <= input(574);
pruneoutput(362) <= input(575);
pruneoutput(363) <= input(576);
pruneoutput(364) <= input(580);
pruneoutput(365) <= input(582);
pruneoutput(366) <= input(583);
pruneoutput(367) <= input(584);
pruneoutput(368) <= input(585);
pruneoutput(369) <= input(587);
pruneoutput(370) <= input(588);
pruneoutput(371) <= input(589);
pruneoutput(372) <= input(590);
pruneoutput(373) <= input(591);
pruneoutput(374) <= input(594);
pruneoutput(375) <= input(595);
pruneoutput(376) <= input(596);
pruneoutput(377) <= input(597);
pruneoutput(378) <= input(598);
pruneoutput(379) <= input(601);
pruneoutput(380) <= input(602);
pruneoutput(381) <= input(603);
pruneoutput(382) <= input(604);
pruneoutput(383) <= input(607);
pruneoutput(384) <= input(608);
pruneoutput(385) <= input(609);
pruneoutput(386) <= input(611);
pruneoutput(387) <= input(612);
pruneoutput(388) <= input(615);
pruneoutput(389) <= input(616);
pruneoutput(390) <= input(619);
pruneoutput(391) <= input(620);
pruneoutput(392) <= input(626);
pruneoutput(393) <= input(628);
pruneoutput(394) <= input(629);
pruneoutput(395) <= input(630);
pruneoutput(396) <= input(631);
pruneoutput(397) <= input(632);
pruneoutput(398) <= input(633);
pruneoutput(399) <= input(634);
pruneoutput(400) <= input(637);
pruneoutput(401) <= input(638);
pruneoutput(402) <= input(639);
pruneoutput(403) <= input(640);
pruneoutput(404) <= input(641);
pruneoutput(405) <= input(642);
pruneoutput(406) <= input(643);
pruneoutput(407) <= input(644);
pruneoutput(408) <= input(645);
pruneoutput(409) <= input(646);
pruneoutput(410) <= input(648);
pruneoutput(411) <= input(649);
pruneoutput(412) <= input(650);
pruneoutput(413) <= input(651);
pruneoutput(414) <= input(652);
pruneoutput(415) <= input(656);
pruneoutput(416) <= input(665);
pruneoutput(417) <= input(667);
pruneoutput(418) <= input(668);
pruneoutput(419) <= input(669);
pruneoutput(420) <= input(670);
pruneoutput(421) <= input(671);
pruneoutput(422) <= input(672);
pruneoutput(423) <= input(674);
pruneoutput(424) <= input(675);
pruneoutput(425) <= input(676);
pruneoutput(426) <= input(677);
pruneoutput(427) <= input(678);
pruneoutput(428) <= input(679);
pruneoutput(429) <= input(680);
pruneoutput(430) <= input(681);
pruneoutput(431) <= input(682);
pruneoutput(432) <= input(683);
pruneoutput(433) <= input(684);
pruneoutput(434) <= input(687);
pruneoutput(435) <= input(688);
pruneoutput(436) <= input(689);
pruneoutput(437) <= input(694);
pruneoutput(438) <= input(695);
pruneoutput(439) <= input(696);
pruneoutput(440) <= input(697);
pruneoutput(441) <= input(698);
pruneoutput(442) <= input(699);
pruneoutput(443) <= input(700);
pruneoutput(444) <= input(701);
pruneoutput(445) <= input(703);
pruneoutput(446) <= input(704);
pruneoutput(447) <= input(706);
pruneoutput(448) <= input(707);
pruneoutput(449) <= input(708);
pruneoutput(450) <= input(710);
pruneoutput(451) <= input(712);
pruneoutput(452) <= input(713);
pruneoutput(453) <= input(716);
pruneoutput(454) <= input(717);
pruneoutput(455) <= input(718);
pruneoutput(456) <= input(719);
pruneoutput(457) <= input(720);
pruneoutput(458) <= input(721);
pruneoutput(459) <= input(723);
pruneoutput(460) <= input(725);
pruneoutput(461) <= input(726);
pruneoutput(462) <= input(727);
pruneoutput(463) <= input(728);
pruneoutput(464) <= input(729);
pruneoutput(465) <= input(730);
pruneoutput(466) <= input(731);
pruneoutput(467) <= input(732);
pruneoutput(468) <= input(734);
pruneoutput(469) <= input(735);
pruneoutput(470) <= input(736);
pruneoutput(471) <= input(737);
pruneoutput(472) <= input(738);
pruneoutput(473) <= input(739);
pruneoutput(474) <= input(740);
pruneoutput(475) <= input(741);
pruneoutput(476) <= input(742);
pruneoutput(477) <= input(743);
pruneoutput(478) <= input(744);
pruneoutput(479) <= input(745);
pruneoutput(480) <= input(751);
pruneoutput(481) <= input(752);
pruneoutput(482) <= input(753);
pruneoutput(483) <= input(754);
pruneoutput(484) <= input(755);
pruneoutput(485) <= input(756);
pruneoutput(486) <= input(757);
pruneoutput(487) <= input(758);
pruneoutput(488) <= input(759);
pruneoutput(489) <= input(760);
pruneoutput(490) <= input(761);
pruneoutput(491) <= input(762);
pruneoutput(492) <= input(763);
pruneoutput(493) <= input(764);
pruneoutput(494) <= input(765);
pruneoutput(495) <= input(766);
pruneoutput(496) <= input(767);
pruneoutput(497) <= input(768);
pruneoutput(498) <= input(769);
pruneoutput(499) <= input(770);
pruneoutput(500) <= input(773);
pruneoutput(501) <= input(774);
pruneoutput(502) <= input(775);
pruneoutput(503) <= input(776);
pruneoutput(504) <= input(777);
pruneoutput(505) <= input(778);
pruneoutput(506) <= input(779);
pruneoutput(507) <= input(780);
pruneoutput(508) <= input(781);
pruneoutput(509) <= input(782);
pruneoutput(510) <= input(783);
pruneoutput(511) <= input(787);
pruneoutput(512) <= input(788);
pruneoutput(513) <= input(789);
pruneoutput(514) <= input(790);
pruneoutput(515) <= input(791);
pruneoutput(516) <= input(792);
pruneoutput(517) <= input(794);
pruneoutput(518) <= input(795);
pruneoutput(519) <= input(796);
pruneoutput(520) <= input(797);
pruneoutput(521) <= input(798);
pruneoutput(522) <= input(799);
pruneoutput(523) <= input(800);
pruneoutput(524) <= input(803);
pruneoutput(525) <= input(804);
pruneoutput(526) <= input(805);
pruneoutput(527) <= input(806);
pruneoutput(528) <= input(807);
pruneoutput(529) <= input(808);
pruneoutput(530) <= input(809);
pruneoutput(531) <= input(810);
pruneoutput(532) <= input(811);
pruneoutput(533) <= input(812);
pruneoutput(534) <= input(813);
pruneoutput(535) <= input(814);
pruneoutput(536) <= input(818);
pruneoutput(537) <= input(819);
pruneoutput(538) <= input(820);
pruneoutput(539) <= input(821);
pruneoutput(540) <= input(822);
pruneoutput(541) <= input(823);
pruneoutput(542) <= input(824);
pruneoutput(543) <= input(825);
pruneoutput(544) <= input(826);
pruneoutput(545) <= input(830);
pruneoutput(546) <= input(831);
pruneoutput(547) <= input(832);
pruneoutput(548) <= input(833);
pruneoutput(549) <= input(834);
pruneoutput(550) <= input(835);
pruneoutput(551) <= input(836);
pruneoutput(552) <= input(841);
pruneoutput(553) <= input(845);
pruneoutput(554) <= input(846);
pruneoutput(555) <= input(847);
pruneoutput(556) <= input(852);
pruneoutput(557) <= input(853);
pruneoutput(558) <= input(854);
pruneoutput(559) <= input(855);
pruneoutput(560) <= input(856);
pruneoutput(561) <= input(857);
pruneoutput(562) <= input(858);
pruneoutput(563) <= input(864);
pruneoutput(564) <= input(865);
pruneoutput(565) <= input(867);
pruneoutput(566) <= input(878);
pruneoutput(567) <= input(879);
pruneoutput(568) <= input(883);
pruneoutput(569) <= input(884);
pruneoutput(570) <= input(885);
pruneoutput(571) <= input(886);
pruneoutput(572) <= input(887);
pruneoutput(573) <= input(891);
pruneoutput(574) <= input(892);
pruneoutput(575) <= input(894);
pruneoutput(576) <= input(897);
pruneoutput(577) <= input(898);
pruneoutput(578) <= input(899);
pruneoutput(579) <= input(900);
pruneoutput(580) <= input(902);
pruneoutput(581) <= input(903);
pruneoutput(582) <= input(904);
pruneoutput(583) <= input(909);
pruneoutput(584) <= input(911);
pruneoutput(585) <= input(912);
pruneoutput(586) <= input(913);
pruneoutput(587) <= input(914);
pruneoutput(588) <= input(915);
pruneoutput(589) <= input(916);
pruneoutput(590) <= input(917);
pruneoutput(591) <= input(918);
pruneoutput(592) <= input(921);
pruneoutput(593) <= input(922);
pruneoutput(594) <= input(923);
pruneoutput(595) <= input(924);
pruneoutput(596) <= input(925);
pruneoutput(597) <= input(926);
pruneoutput(598) <= input(927);
pruneoutput(599) <= input(928);
pruneoutput(600) <= input(929);
pruneoutput(601) <= input(930);
pruneoutput(602) <= input(931);
pruneoutput(603) <= input(932);
pruneoutput(604) <= input(933);
pruneoutput(605) <= input(934);
pruneoutput(606) <= input(935);
pruneoutput(607) <= input(936);
pruneoutput(608) <= input(937);
pruneoutput(609) <= input(938);
pruneoutput(610) <= input(939);
pruneoutput(611) <= input(946);
pruneoutput(612) <= input(948);
pruneoutput(613) <= input(949);
pruneoutput(614) <= input(950);
pruneoutput(615) <= input(951);
pruneoutput(616) <= input(952);
pruneoutput(617) <= input(953);
pruneoutput(618) <= input(954);
pruneoutput(619) <= input(955);
pruneoutput(620) <= input(956);
pruneoutput(621) <= input(957);
pruneoutput(622) <= input(958);
pruneoutput(623) <= input(960);
pruneoutput(624) <= input(961);
pruneoutput(625) <= input(962);
pruneoutput(626) <= input(970);
pruneoutput(627) <= input(973);
pruneoutput(628) <= input(974);
pruneoutput(629) <= input(975);
pruneoutput(630) <= input(976);
pruneoutput(631) <= input(977);
pruneoutput(632) <= input(978);
pruneoutput(633) <= input(979);
pruneoutput(634) <= input(983);
pruneoutput(635) <= input(984);
pruneoutput(636) <= input(985);
pruneoutput(637) <= input(986);
pruneoutput(638) <= input(988);
pruneoutput(639) <= input(989);
pruneoutput(640) <= input(999);

END ARCHITECTURE behavioral;