LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY BasedVectorLFSR IS
	GENERIC ( n	: INTEGER	:= 2000			    -- number of bits
				);	 
	PORT (
		clk, rst, update	: IN STD_LOGIC; 
		congigSignitureIn , congigInitialvaluesIn : IN STD_LOGIC_VECTOR (n-1 DOWNTO 0 );
		dout				: OUT  STD_LOGIC_VECTOR (n-1 DOWNTO 0 )
	);
END ENTITY BasedVectorLFSR;

ARCHITECTURE behavioral OF BasedVectorLFSR IS

COMPONENT  regOne IS
	GENERIC (init : STD_LOGIC := '1');   -- initial value
	PORT (
		clk 				: IN  STD_LOGIC;
		regUpdate, regrst 	: IN  STD_LOGIC;
		din        			: IN  STD_LOGIC;
		dout        		: OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL interValIn : STD_LOGIC_VECTOR (n-1 DOWNTO 0);
SIGNAL interValOut : STD_LOGIC_VECTOR (n-1 DOWNTO 0);
SIGNAL interValOutR : STD_LOGIC_VECTOR (0 TO n-1);
CONSTANT congigSigniture : STD_LOGIC_VECTOR (n-1 DOWNTO 0) :=    "1100011001101000001010100111100110101010000110110101010000010010111010000000001001101011000011111100100010011111111110101100010101110101000011101111111101101100111011000001001011111011100000110101001011101000101001011110011000111101001100100100011100101001000000001011010101000110001100101001001011101101110110111010101010101001100001110011010001001110010010010111010000000010010111011110101010010111101101010110100000001101101011011011000001011000010111110111010010111000000011110001010001110101110010001011010010000010000010000010001001001001110101100111011010010110000011011000101010100110000101101011011101111000011001000110101110101011010010111000101010010000100101100100101000010000110100000100111001110111110001111100001110101011100001100111101000000110100010011110001001111000010001001011100010111010110010001000001000001001111000111001010110011111001010100101001101011000111001010010011100100101011100111000001100100101000111011110110100010011011000100111000000110000101011110111010000001011"; --"1010101011000011001011001000001001000110100100000010011011000001110101100010000001000111100011101100011001100110100010101100010001011111010110000011000010111011110110101000110101100100110110100001010010111100101010101000111011111101101111011111001111001010110000010110100001111110011100100000000110110110000000011011010111101011100110101100010100100011010011000001010111000000010001101101101011010110110011110000010000110110010110100011111001011110011010011101011010111100011001010111011111110101100110001110000011111111110110001011001111111110010101010010011101000011100111101011011000110101010101100000100001101010101000111111001001111101010000110001110110001010111000101100101010011110010101100010011011011111111100100111100010011100101010010000001100111011100101101011100010111001000110101111110111111010001000100101100011100010001011001100110111011010101010000010100000000101001000110011011011011100010011011001001011100000000000000001000010010101100101110110001001101010101101010001110000001100";

CONSTANT congigInitialvalues : STD_LOGIC_VECTOR (n-1 DOWNTO 0) := "1100011111100001110000010001110000100000101101000111010010010010110001011101100001100010001111100001111110000011110110000111100001011110111110010011110011100101101010100110001010100101110100111001101100011100110111010000010111011111011101001001111001111110001000010011000000111101100111101001111101111010101010001001000111111110101001011000101010010101011010110100000011110110000111100100110101101111101100110010011010001101010100011011001000011000100100010110110000000010000001000100101111111000101001101000000101111010100100011110001011001101110000011011001110011010110101101111010100010011100010010000000101010001011100101000101010010000110110000000000110010110100011000010111010010011011001101001100000100101001000100000100010000000111011110110111101000110001101001010110100011100111111001110110001100000101000100111101001111101011000100000010100100001110000110100011111011100010010101001100101010110101011011011000010010001101100001011011100110100011110110000001001100011111100111100110111111010";--"1111000000100110110100000110111010000101111100010011000110000110000100100100100010111110100100111000000001010111001001001000111010011010000001011010010100111000100010110111010111110010000101010100011101011111011100001011010100011100110110100001101100111100101111001001100100000011110111000110111000010001111100011110001110001010001011011011000000001010000001000001000011100010110011111101111000000010000111110001101011110111101010101010001110110110100100101011011011011110000111110110011000100110111010000011101100111010000010101011010111001011110110100000101100101111110011010011010010111000100100101100101101010001001110100010100001011100010111110010110011101000111110110001100100011100001110110000101111110011100100011011011101101110010101000101010100101011110011100100111100010011011100100101001010000110000101011100001110011111100011000011101010100001011010100101011110000100010001101001000000001011010001001001001000111010110101000010101011111110000010001010100111111100100011000110110101100110";

BEGIN

	regArr : FOR i IN 1 TO n-1 GENERATE
		Ireg : regOne 
			GENERIC map(congigInitialvalues(i))
			PORT map(clk,  update, rst, 
			interValIn(i), 	interValOut(i) 
					 );   
	END GENERATE regArr;
	xorchain : FOR i IN 1 TO n-1 GENERATE
	xorchain1: IF (congigSigniture(i) = '1') GENERATE
			interValIn(i) <= interValOut(i-1) XOR  interValOut(n-1);
		END GENERATE xorchain1;
	xorchain2: IF (congigSigniture(i) = '0') GENERATE
			interValIn(i) <= interValOut(i-1);
		END GENERATE xorchain2;
	END GENERATE xorchain;
	interValIn(0) <= interValOut(n-1);
	reg0 : regOne 
			GENERIC map(congigInitialvalues(0))
			PORT map(clk,  update, rst, 
			interValIn(0), 	interValOut(0) 
					 ); 
	--interValOutR <= interValOut;
	dout <= interValOut;--(0 TO n-1);

END ARCHITECTURE behavioral;