LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY BasedVectorLFSR IS
	GENERIC ( n	: INTEGER	:= 2000;			    -- number of bits
			  s	: INTEGER	:= 8;   		    -- signiture in decimal 
			  i	: INTEGER	:= 8    		    -- initialvalues in decimal 
				);	 
	PORT (
		clk, rst, update	: IN STD_LOGIC; 
		dout				: OUT  STD_LOGIC_VECTOR (n-1 DOWNTO 0 )
	);
END ENTITY BasedVectorLFSR;

ARCHITECTURE behavioral OF BasedVectorLFSR IS

COMPONENT  regOne IS
	GENERIC (init : STD_LOGIC := '1');   -- initial value
	PORT (
		clk 				: IN  STD_LOGIC;
		regUpdate, regrst 	: IN  STD_LOGIC;
		din        			: IN  STD_LOGIC;
		dout        		: OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL interValIn : STD_LOGIC_VECTOR (n-1 DOWNTO 0);
SIGNAL interValOut : STD_LOGIC_VECTOR (n-1 DOWNTO 0);
SIGNAL interValOutR : STD_LOGIC_VECTOR (0 TO n-1);
CONSTANT congigSigniture : STD_LOGIC_VECTOR (n-1 DOWNTO 0) :=    "1110001100011110011110001111110000111111001101101011011001001000111100001001100000110001101010101111001101001111000111010100100100110000110010111110010010010111000010001000111010010011110000001101100001110101100000111110000011100000011111110010011100110100011010000100010000111000000111101001001001111001000101001000101101111110001000101010000010010010100011010101011001110011100101110000010110001101110100110001111110111111111010000110101110110110101110110000001110101101101111011011011011100000000110001011010011001010111011001111000011101100011010000111110010111111011001001100000110000000000001111010010110100001000011011010001011010000011110000000100011000000011011000011011010111100010011111001101001110100111111001111101001011100100010010010010111000110001000101100101101001100101101010001101001010100110000000110101100110111100010100010001000101100010100011000001110101000100000011000001110011101111001001101000011101101100001110110111101010111110111011000000111001100010110101000010011010001";

CONSTANT congigInitialvalues : STD_LOGIC_VECTOR (n-1 DOWNTO 0):= "0111100100110101101001000101100010111111111100100100100100001011101001100010000111111010001001111011110110100000101110111101101000110010011001010011101010100110010011111011011001111000110101111011101111100101101001000101110011101100101000110100001010000011100100010110100100100010111001101001000111001000000100111011000010001100101011001000101011011000111011011000001110000001100010110110000100001011100011001110110101100111011011100001001100011001011010000100000001110100000111100010100110010011101110101111111100000101110101111111010010010101011011001111100110001011010101110111011110101100111111010010000111010001011010001000101011101000001111001101101011011000001111010110000110010001110001010010000111000000110100001100001111110001111010001100110010111100011010000010011101000010000011111010100110110110000100011110100011001000000100100000001111011110100100111110100111010110100011011011001010110101100100111011101111001011101100010111100100000101010100001110011001000101001111110111011001010001";
---- 0111100100110101101001000101100010111111111100100100100100001011101001100010000111111010001001111011110110100000101110111101101000110010011001010011101010100110010011111011011001111000110101111011101111100101101001000101110011101100101000110100001010000011100100010110100100100010111001101001000111001000000100111011000010001100101011001000101011011000111011011000001110000001100010110110000100001011100011001110110101100111011011100001001100011001011010000100000001110100000111100010100110010011101110101111111100000101110101111111010010010101011011001111100110001011010101110111011110101100111111010010000111010001011010001000101011101000001111001101101011011000001111010110000110010001110001010010000111000000110100001100001111110001111010001100110010111100011010000010011101000010000011111010100110110110000100011110100011001000000100100000001111011110100100111110100111010110100011011011001010110101100100111011101111001011101100010111100100000101010100001110011001000101001111110111011001010001
----- orgINIT 1110001100011110011110001111110000111111001101101011011001001000111100001001100000110001101010101111001101001111000111010100100100110000110010111110010010010111000010001000111010010011110000001101100001110101100000111110000011100000011111110010011100110100011010000100010000111000000111101001001001111001000101001000101101111110001000101010000010010010100011010101011001110011100101110000010110001101110100110001111110111111111010000110101110110110101110110000001110101101101111011011011011100000000110001011010011001010111011001111000011101100011010000111110010111111011001001100000110000000000001111010010110100001000011011010001011010000011110000000100011000000011011000011011010111100010011111001101001110100111111001111101001011100100010010010010111000110001000101100101101001100101101010001101001010100110000000110101100110111100010100010001000101100010100011000001110101000100000011000001110011101111001001101000011101101100001110110111101010111110111011000000111001100010110101000010011010001
BEGIN


	regArr : FOR i IN 1 TO n-1 GENERATE
		Ireg : regOne 
			GENERIC map(congigInitialvalues(i))
			PORT map(clk,  update, rst, 
			interValIn(i), 	interValOut(i) 
					 );   
	END GENERATE regArr;
	xorchain : FOR i IN 1 TO n-1 GENERATE
	xorchain1: IF (congigSigniture(i) = '1') GENERATE
			interValIn(i) <= interValOut(i-1) XOR  interValOut(n-1);
		END GENERATE xorchain1;
	xorchain2: IF (congigSigniture(i) = '0') GENERATE
			interValIn(i) <= interValOut(i-1);
		END GENERATE xorchain2;
	END GENERATE xorchain;
	interValIn(0) <= interValOut(n-1);
	reg0 : regOne 
			GENERIC map(congigInitialvalues(0))
			PORT map(clk,  update, rst, 
			interValIn(0), 	interValOut(0) 
					 ); 
	--interValOutR <= interValOut;
	dout <= interValOut;--(0 TO n-1);

END ARCHITECTURE behavioral;
-------------------------------------------------------------------------------
