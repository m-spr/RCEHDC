LIBRARY IEEE; 
USE IEEE.STD_LOGIC_1164.ALL; 
USE IEEE.NUMERIC_STD.ALL; 
  
ENTITY connector IS 
	PORT ( 
		input         : IN  STD_LOGIC_VECTOR (1099 DOWNTO 0); 
		pruneoutput        : OUT  STD_LOGIC_VECTOR (679 DOWNTO 0)      
	);
END ENTITY connector;

ARCHITECTURE behavioral OF connector  IS
BEGIN
pruneoutput(0) <= input(3);
pruneoutput(1) <= input(4);
pruneoutput(2) <= input(5);
pruneoutput(3) <= input(7);
pruneoutput(4) <= input(9);
pruneoutput(5) <= input(12);
pruneoutput(6) <= input(13);
pruneoutput(7) <= input(14);
pruneoutput(8) <= input(15);
pruneoutput(9) <= input(16);
pruneoutput(10) <= input(17);
pruneoutput(11) <= input(18);
pruneoutput(12) <= input(22);
pruneoutput(13) <= input(23);
pruneoutput(14) <= input(25);
pruneoutput(15) <= input(30);
pruneoutput(16) <= input(31);
pruneoutput(17) <= input(34);
pruneoutput(18) <= input(35);
pruneoutput(19) <= input(36);
pruneoutput(20) <= input(39);
pruneoutput(21) <= input(40);
pruneoutput(22) <= input(41);
pruneoutput(23) <= input(42);
pruneoutput(24) <= input(48);
pruneoutput(25) <= input(49);
pruneoutput(26) <= input(50);
pruneoutput(27) <= input(54);
pruneoutput(28) <= input(55);
pruneoutput(29) <= input(56);
pruneoutput(30) <= input(57);
pruneoutput(31) <= input(60);
pruneoutput(32) <= input(61);
pruneoutput(33) <= input(62);
pruneoutput(34) <= input(63);
pruneoutput(35) <= input(76);
pruneoutput(36) <= input(77);
pruneoutput(37) <= input(78);
pruneoutput(38) <= input(79);
pruneoutput(39) <= input(80);
pruneoutput(40) <= input(81);
pruneoutput(41) <= input(82);
pruneoutput(42) <= input(83);
pruneoutput(43) <= input(87);
pruneoutput(44) <= input(88);
pruneoutput(45) <= input(91);
pruneoutput(46) <= input(92);
pruneoutput(47) <= input(93);
pruneoutput(48) <= input(94);
pruneoutput(49) <= input(95);
pruneoutput(50) <= input(96);
pruneoutput(51) <= input(98);
pruneoutput(52) <= input(99);
pruneoutput(53) <= input(100);
pruneoutput(54) <= input(104);
pruneoutput(55) <= input(105);
pruneoutput(56) <= input(106);
pruneoutput(57) <= input(107);
pruneoutput(58) <= input(108);
pruneoutput(59) <= input(109);
pruneoutput(60) <= input(110);
pruneoutput(61) <= input(111);
pruneoutput(62) <= input(112);
pruneoutput(63) <= input(113);
pruneoutput(64) <= input(114);
pruneoutput(65) <= input(120);
pruneoutput(66) <= input(121);
pruneoutput(67) <= input(123);
pruneoutput(68) <= input(124);
pruneoutput(69) <= input(125);
pruneoutput(70) <= input(126);
pruneoutput(71) <= input(127);
pruneoutput(72) <= input(128);
pruneoutput(73) <= input(129);
pruneoutput(74) <= input(130);
pruneoutput(75) <= input(131);
pruneoutput(76) <= input(136);
pruneoutput(77) <= input(137);
pruneoutput(78) <= input(138);
pruneoutput(79) <= input(139);
pruneoutput(80) <= input(140);
pruneoutput(81) <= input(141);
pruneoutput(82) <= input(142);
pruneoutput(83) <= input(143);
pruneoutput(84) <= input(144);
pruneoutput(85) <= input(145);
pruneoutput(86) <= input(146);
pruneoutput(87) <= input(147);
pruneoutput(88) <= input(148);
pruneoutput(89) <= input(149);
pruneoutput(90) <= input(150);
pruneoutput(91) <= input(151);
pruneoutput(92) <= input(153);
pruneoutput(93) <= input(154);
pruneoutput(94) <= input(156);
pruneoutput(95) <= input(157);
pruneoutput(96) <= input(160);
pruneoutput(97) <= input(161);
pruneoutput(98) <= input(162);
pruneoutput(99) <= input(166);
pruneoutput(100) <= input(167);
pruneoutput(101) <= input(169);
pruneoutput(102) <= input(171);
pruneoutput(103) <= input(174);
pruneoutput(104) <= input(175);
pruneoutput(105) <= input(176);
pruneoutput(106) <= input(178);
pruneoutput(107) <= input(185);
pruneoutput(108) <= input(186);
pruneoutput(109) <= input(187);
pruneoutput(110) <= input(188);
pruneoutput(111) <= input(189);
pruneoutput(112) <= input(190);
pruneoutput(113) <= input(191);
pruneoutput(114) <= input(192);
pruneoutput(115) <= input(193);
pruneoutput(116) <= input(198);
pruneoutput(117) <= input(199);
pruneoutput(118) <= input(203);
pruneoutput(119) <= input(204);
pruneoutput(120) <= input(205);
pruneoutput(121) <= input(206);
pruneoutput(122) <= input(209);
pruneoutput(123) <= input(212);
pruneoutput(124) <= input(214);
pruneoutput(125) <= input(215);
pruneoutput(126) <= input(216);
pruneoutput(127) <= input(217);
pruneoutput(128) <= input(218);
pruneoutput(129) <= input(219);
pruneoutput(130) <= input(220);
pruneoutput(131) <= input(225);
pruneoutput(132) <= input(226);
pruneoutput(133) <= input(227);
pruneoutput(134) <= input(232);
pruneoutput(135) <= input(233);
pruneoutput(136) <= input(236);
pruneoutput(137) <= input(237);
pruneoutput(138) <= input(238);
pruneoutput(139) <= input(239);
pruneoutput(140) <= input(240);
pruneoutput(141) <= input(241);
pruneoutput(142) <= input(242);
pruneoutput(143) <= input(245);
pruneoutput(144) <= input(246);
pruneoutput(145) <= input(247);
pruneoutput(146) <= input(248);
pruneoutput(147) <= input(249);
pruneoutput(148) <= input(250);
pruneoutput(149) <= input(251);
pruneoutput(150) <= input(253);
pruneoutput(151) <= input(254);
pruneoutput(152) <= input(255);
pruneoutput(153) <= input(256);
pruneoutput(154) <= input(257);
pruneoutput(155) <= input(258);
pruneoutput(156) <= input(261);
pruneoutput(157) <= input(262);
pruneoutput(158) <= input(263);
pruneoutput(159) <= input(265);
pruneoutput(160) <= input(266);
pruneoutput(161) <= input(267);
pruneoutput(162) <= input(275);
pruneoutput(163) <= input(276);
pruneoutput(164) <= input(277);
pruneoutput(165) <= input(278);
pruneoutput(166) <= input(280);
pruneoutput(167) <= input(281);
pruneoutput(168) <= input(282);
pruneoutput(169) <= input(283);
pruneoutput(170) <= input(284);
pruneoutput(171) <= input(288);
pruneoutput(172) <= input(289);
pruneoutput(173) <= input(290);
pruneoutput(174) <= input(291);
pruneoutput(175) <= input(292);
pruneoutput(176) <= input(294);
pruneoutput(177) <= input(296);
pruneoutput(178) <= input(298);
pruneoutput(179) <= input(306);
pruneoutput(180) <= input(307);
pruneoutput(181) <= input(308);
pruneoutput(182) <= input(309);
pruneoutput(183) <= input(312);
pruneoutput(184) <= input(313);
pruneoutput(185) <= input(314);
pruneoutput(186) <= input(321);
pruneoutput(187) <= input(322);
pruneoutput(188) <= input(326);
pruneoutput(189) <= input(330);
pruneoutput(190) <= input(331);
pruneoutput(191) <= input(332);
pruneoutput(192) <= input(333);
pruneoutput(193) <= input(334);
pruneoutput(194) <= input(335);
pruneoutput(195) <= input(336);
pruneoutput(196) <= input(337);
pruneoutput(197) <= input(341);
pruneoutput(198) <= input(342);
pruneoutput(199) <= input(343);
pruneoutput(200) <= input(344);
pruneoutput(201) <= input(345);
pruneoutput(202) <= input(346);
pruneoutput(203) <= input(347);
pruneoutput(204) <= input(349);
pruneoutput(205) <= input(350);
pruneoutput(206) <= input(351);
pruneoutput(207) <= input(353);
pruneoutput(208) <= input(354);
pruneoutput(209) <= input(355);
pruneoutput(210) <= input(356);
pruneoutput(211) <= input(359);
pruneoutput(212) <= input(360);
pruneoutput(213) <= input(361);
pruneoutput(214) <= input(362);
pruneoutput(215) <= input(363);
pruneoutput(216) <= input(364);
pruneoutput(217) <= input(365);
pruneoutput(218) <= input(366);
pruneoutput(219) <= input(367);
pruneoutput(220) <= input(368);
pruneoutput(221) <= input(369);
pruneoutput(222) <= input(370);
pruneoutput(223) <= input(371);
pruneoutput(224) <= input(372);
pruneoutput(225) <= input(375);
pruneoutput(226) <= input(376);
pruneoutput(227) <= input(378);
pruneoutput(228) <= input(379);
pruneoutput(229) <= input(384);
pruneoutput(230) <= input(389);
pruneoutput(231) <= input(390);
pruneoutput(232) <= input(391);
pruneoutput(233) <= input(396);
pruneoutput(234) <= input(397);
pruneoutput(235) <= input(398);
pruneoutput(236) <= input(399);
pruneoutput(237) <= input(402);
pruneoutput(238) <= input(403);
pruneoutput(239) <= input(404);
pruneoutput(240) <= input(406);
pruneoutput(241) <= input(407);
pruneoutput(242) <= input(413);
pruneoutput(243) <= input(414);
pruneoutput(244) <= input(415);
pruneoutput(245) <= input(417);
pruneoutput(246) <= input(418);
pruneoutput(247) <= input(419);
pruneoutput(248) <= input(420);
pruneoutput(249) <= input(421);
pruneoutput(250) <= input(422);
pruneoutput(251) <= input(423);
pruneoutput(252) <= input(424);
pruneoutput(253) <= input(428);
pruneoutput(254) <= input(429);
pruneoutput(255) <= input(430);
pruneoutput(256) <= input(431);
pruneoutput(257) <= input(435);
pruneoutput(258) <= input(436);
pruneoutput(259) <= input(437);
pruneoutput(260) <= input(439);
pruneoutput(261) <= input(440);
pruneoutput(262) <= input(441);
pruneoutput(263) <= input(442);
pruneoutput(264) <= input(443);
pruneoutput(265) <= input(444);
pruneoutput(266) <= input(446);
pruneoutput(267) <= input(447);
pruneoutput(268) <= input(448);
pruneoutput(269) <= input(449);
pruneoutput(270) <= input(450);
pruneoutput(271) <= input(451);
pruneoutput(272) <= input(453);
pruneoutput(273) <= input(454);
pruneoutput(274) <= input(455);
pruneoutput(275) <= input(456);
pruneoutput(276) <= input(457);
pruneoutput(277) <= input(458);
pruneoutput(278) <= input(459);
pruneoutput(279) <= input(460);
pruneoutput(280) <= input(461);
pruneoutput(281) <= input(466);
pruneoutput(282) <= input(469);
pruneoutput(283) <= input(476);
pruneoutput(284) <= input(478);
pruneoutput(285) <= input(479);
pruneoutput(286) <= input(480);
pruneoutput(287) <= input(481);
pruneoutput(288) <= input(482);
pruneoutput(289) <= input(483);
pruneoutput(290) <= input(484);
pruneoutput(291) <= input(485);
pruneoutput(292) <= input(487);
pruneoutput(293) <= input(488);
pruneoutput(294) <= input(489);
pruneoutput(295) <= input(490);
pruneoutput(296) <= input(491);
pruneoutput(297) <= input(492);
pruneoutput(298) <= input(493);
pruneoutput(299) <= input(494);
pruneoutput(300) <= input(496);
pruneoutput(301) <= input(497);
pruneoutput(302) <= input(498);
pruneoutput(303) <= input(499);
pruneoutput(304) <= input(500);
pruneoutput(305) <= input(501);
pruneoutput(306) <= input(503);
pruneoutput(307) <= input(510);
pruneoutput(308) <= input(511);
pruneoutput(309) <= input(515);
pruneoutput(310) <= input(520);
pruneoutput(311) <= input(524);
pruneoutput(312) <= input(525);
pruneoutput(313) <= input(529);
pruneoutput(314) <= input(530);
pruneoutput(315) <= input(531);
pruneoutput(316) <= input(532);
pruneoutput(317) <= input(533);
pruneoutput(318) <= input(534);
pruneoutput(319) <= input(535);
pruneoutput(320) <= input(536);
pruneoutput(321) <= input(537);
pruneoutput(322) <= input(538);
pruneoutput(323) <= input(539);
pruneoutput(324) <= input(540);
pruneoutput(325) <= input(542);
pruneoutput(326) <= input(543);
pruneoutput(327) <= input(544);
pruneoutput(328) <= input(545);
pruneoutput(329) <= input(546);
pruneoutput(330) <= input(547);
pruneoutput(331) <= input(551);
pruneoutput(332) <= input(552);
pruneoutput(333) <= input(553);
pruneoutput(334) <= input(554);
pruneoutput(335) <= input(557);
pruneoutput(336) <= input(558);
pruneoutput(337) <= input(561);
pruneoutput(338) <= input(562);
pruneoutput(339) <= input(566);
pruneoutput(340) <= input(569);
pruneoutput(341) <= input(570);
pruneoutput(342) <= input(572);
pruneoutput(343) <= input(573);
pruneoutput(344) <= input(574);
pruneoutput(345) <= input(580);
pruneoutput(346) <= input(585);
pruneoutput(347) <= input(586);
pruneoutput(348) <= input(588);
pruneoutput(349) <= input(589);
pruneoutput(350) <= input(590);
pruneoutput(351) <= input(591);
pruneoutput(352) <= input(593);
pruneoutput(353) <= input(594);
pruneoutput(354) <= input(595);
pruneoutput(355) <= input(596);
pruneoutput(356) <= input(597);
pruneoutput(357) <= input(598);
pruneoutput(358) <= input(599);
pruneoutput(359) <= input(600);
pruneoutput(360) <= input(601);
pruneoutput(361) <= input(602);
pruneoutput(362) <= input(603);
pruneoutput(363) <= input(604);
pruneoutput(364) <= input(605);
pruneoutput(365) <= input(606);
pruneoutput(366) <= input(607);
pruneoutput(367) <= input(608);
pruneoutput(368) <= input(609);
pruneoutput(369) <= input(610);
pruneoutput(370) <= input(611);
pruneoutput(371) <= input(612);
pruneoutput(372) <= input(614);
pruneoutput(373) <= input(619);
pruneoutput(374) <= input(620);
pruneoutput(375) <= input(621);
pruneoutput(376) <= input(622);
pruneoutput(377) <= input(623);
pruneoutput(378) <= input(624);
pruneoutput(379) <= input(625);
pruneoutput(380) <= input(626);
pruneoutput(381) <= input(627);
pruneoutput(382) <= input(628);
pruneoutput(383) <= input(629);
pruneoutput(384) <= input(630);
pruneoutput(385) <= input(631);
pruneoutput(386) <= input(632);
pruneoutput(387) <= input(633);
pruneoutput(388) <= input(634);
pruneoutput(389) <= input(635);
pruneoutput(390) <= input(636);
pruneoutput(391) <= input(637);
pruneoutput(392) <= input(638);
pruneoutput(393) <= input(639);
pruneoutput(394) <= input(640);
pruneoutput(395) <= input(641);
pruneoutput(396) <= input(642);
pruneoutput(397) <= input(643);
pruneoutput(398) <= input(644);
pruneoutput(399) <= input(647);
pruneoutput(400) <= input(648);
pruneoutput(401) <= input(649);
pruneoutput(402) <= input(651);
pruneoutput(403) <= input(652);
pruneoutput(404) <= input(656);
pruneoutput(405) <= input(657);
pruneoutput(406) <= input(658);
pruneoutput(407) <= input(659);
pruneoutput(408) <= input(660);
pruneoutput(409) <= input(661);
pruneoutput(410) <= input(662);
pruneoutput(411) <= input(667);
pruneoutput(412) <= input(671);
pruneoutput(413) <= input(672);
pruneoutput(414) <= input(673);
pruneoutput(415) <= input(674);
pruneoutput(416) <= input(675);
pruneoutput(417) <= input(676);
pruneoutput(418) <= input(677);
pruneoutput(419) <= input(678);
pruneoutput(420) <= input(681);
pruneoutput(421) <= input(682);
pruneoutput(422) <= input(683);
pruneoutput(423) <= input(684);
pruneoutput(424) <= input(685);
pruneoutput(425) <= input(686);
pruneoutput(426) <= input(687);
pruneoutput(427) <= input(688);
pruneoutput(428) <= input(689);
pruneoutput(429) <= input(690);
pruneoutput(430) <= input(691);
pruneoutput(431) <= input(692);
pruneoutput(432) <= input(693);
pruneoutput(433) <= input(695);
pruneoutput(434) <= input(696);
pruneoutput(435) <= input(697);
pruneoutput(436) <= input(698);
pruneoutput(437) <= input(705);
pruneoutput(438) <= input(706);
pruneoutput(439) <= input(707);
pruneoutput(440) <= input(708);
pruneoutput(441) <= input(709);
pruneoutput(442) <= input(710);
pruneoutput(443) <= input(711);
pruneoutput(444) <= input(712);
pruneoutput(445) <= input(713);
pruneoutput(446) <= input(714);
pruneoutput(447) <= input(715);
pruneoutput(448) <= input(716);
pruneoutput(449) <= input(720);
pruneoutput(450) <= input(721);
pruneoutput(451) <= input(726);
pruneoutput(452) <= input(731);
pruneoutput(453) <= input(732);
pruneoutput(454) <= input(733);
pruneoutput(455) <= input(737);
pruneoutput(456) <= input(740);
pruneoutput(457) <= input(742);
pruneoutput(458) <= input(743);
pruneoutput(459) <= input(747);
pruneoutput(460) <= input(748);
pruneoutput(461) <= input(750);
pruneoutput(462) <= input(751);
pruneoutput(463) <= input(752);
pruneoutput(464) <= input(753);
pruneoutput(465) <= input(756);
pruneoutput(466) <= input(757);
pruneoutput(467) <= input(758);
pruneoutput(468) <= input(759);
pruneoutput(469) <= input(760);
pruneoutput(470) <= input(761);
pruneoutput(471) <= input(762);
pruneoutput(472) <= input(766);
pruneoutput(473) <= input(767);
pruneoutput(474) <= input(776);
pruneoutput(475) <= input(777);
pruneoutput(476) <= input(778);
pruneoutput(477) <= input(780);
pruneoutput(478) <= input(781);
pruneoutput(479) <= input(782);
pruneoutput(480) <= input(783);
pruneoutput(481) <= input(785);
pruneoutput(482) <= input(786);
pruneoutput(483) <= input(787);
pruneoutput(484) <= input(788);
pruneoutput(485) <= input(789);
pruneoutput(486) <= input(790);
pruneoutput(487) <= input(792);
pruneoutput(488) <= input(793);
pruneoutput(489) <= input(794);
pruneoutput(490) <= input(795);
pruneoutput(491) <= input(796);
pruneoutput(492) <= input(797);
pruneoutput(493) <= input(798);
pruneoutput(494) <= input(804);
pruneoutput(495) <= input(805);
pruneoutput(496) <= input(806);
pruneoutput(497) <= input(807);
pruneoutput(498) <= input(810);
pruneoutput(499) <= input(811);
pruneoutput(500) <= input(812);
pruneoutput(501) <= input(816);
pruneoutput(502) <= input(817);
pruneoutput(503) <= input(818);
pruneoutput(504) <= input(819);
pruneoutput(505) <= input(820);
pruneoutput(506) <= input(821);
pruneoutput(507) <= input(823);
pruneoutput(508) <= input(824);
pruneoutput(509) <= input(825);
pruneoutput(510) <= input(826);
pruneoutput(511) <= input(827);
pruneoutput(512) <= input(828);
pruneoutput(513) <= input(829);
pruneoutput(514) <= input(833);
pruneoutput(515) <= input(834);
pruneoutput(516) <= input(835);
pruneoutput(517) <= input(842);
pruneoutput(518) <= input(843);
pruneoutput(519) <= input(844);
pruneoutput(520) <= input(845);
pruneoutput(521) <= input(848);
pruneoutput(522) <= input(849);
pruneoutput(523) <= input(854);
pruneoutput(524) <= input(855);
pruneoutput(525) <= input(856);
pruneoutput(526) <= input(857);
pruneoutput(527) <= input(858);
pruneoutput(528) <= input(859);
pruneoutput(529) <= input(860);
pruneoutput(530) <= input(861);
pruneoutput(531) <= input(863);
pruneoutput(532) <= input(864);
pruneoutput(533) <= input(865);
pruneoutput(534) <= input(866);
pruneoutput(535) <= input(867);
pruneoutput(536) <= input(868);
pruneoutput(537) <= input(869);
pruneoutput(538) <= input(871);
pruneoutput(539) <= input(875);
pruneoutput(540) <= input(876);
pruneoutput(541) <= input(877);
pruneoutput(542) <= input(878);
pruneoutput(543) <= input(879);
pruneoutput(544) <= input(880);
pruneoutput(545) <= input(881);
pruneoutput(546) <= input(883);
pruneoutput(547) <= input(884);
pruneoutput(548) <= input(885);
pruneoutput(549) <= input(886);
pruneoutput(550) <= input(888);
pruneoutput(551) <= input(889);
pruneoutput(552) <= input(890);
pruneoutput(553) <= input(891);
pruneoutput(554) <= input(892);
pruneoutput(555) <= input(893);
pruneoutput(556) <= input(894);
pruneoutput(557) <= input(895);
pruneoutput(558) <= input(896);
pruneoutput(559) <= input(897);
pruneoutput(560) <= input(898);
pruneoutput(561) <= input(900);
pruneoutput(562) <= input(901);
pruneoutput(563) <= input(902);
pruneoutput(564) <= input(903);
pruneoutput(565) <= input(904);
pruneoutput(566) <= input(905);
pruneoutput(567) <= input(906);
pruneoutput(568) <= input(910);
pruneoutput(569) <= input(911);
pruneoutput(570) <= input(912);
pruneoutput(571) <= input(913);
pruneoutput(572) <= input(914);
pruneoutput(573) <= input(915);
pruneoutput(574) <= input(916);
pruneoutput(575) <= input(919);
pruneoutput(576) <= input(923);
pruneoutput(577) <= input(924);
pruneoutput(578) <= input(926);
pruneoutput(579) <= input(927);
pruneoutput(580) <= input(928);
pruneoutput(581) <= input(933);
pruneoutput(582) <= input(934);
pruneoutput(583) <= input(935);
pruneoutput(584) <= input(936);
pruneoutput(585) <= input(938);
pruneoutput(586) <= input(939);
pruneoutput(587) <= input(940);
pruneoutput(588) <= input(941);
pruneoutput(589) <= input(947);
pruneoutput(590) <= input(948);
pruneoutput(591) <= input(949);
pruneoutput(592) <= input(950);
pruneoutput(593) <= input(951);
pruneoutput(594) <= input(952);
pruneoutput(595) <= input(953);
pruneoutput(596) <= input(956);
pruneoutput(597) <= input(960);
pruneoutput(598) <= input(962);
pruneoutput(599) <= input(963);
pruneoutput(600) <= input(964);
pruneoutput(601) <= input(965);
pruneoutput(602) <= input(966);
pruneoutput(603) <= input(967);
pruneoutput(604) <= input(970);
pruneoutput(605) <= input(971);
pruneoutput(606) <= input(974);
pruneoutput(607) <= input(975);
pruneoutput(608) <= input(976);
pruneoutput(609) <= input(977);
pruneoutput(610) <= input(979);
pruneoutput(611) <= input(983);
pruneoutput(612) <= input(984);
pruneoutput(613) <= input(985);
pruneoutput(614) <= input(986);
pruneoutput(615) <= input(987);
pruneoutput(616) <= input(988);
pruneoutput(617) <= input(989);
pruneoutput(618) <= input(991);
pruneoutput(619) <= input(992);
pruneoutput(620) <= input(993);
pruneoutput(621) <= input(994);
pruneoutput(622) <= input(996);
pruneoutput(623) <= input(997);

END ARCHITECTURE behavioral;