-- MIT License

-- Copyright (c) 2024 m-spr

-- Permission is hereby granted, free of charge, to any person obtaining a copy
-- of this software and associated documentation files (the "Software"), to deal
-- in the Software without restriction, including without limitation the rights
-- to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
-- copies of the Software, and to permit persons to whom the Software is
-- furnished to do so, subject to the following conditions:

-- The above copyright notice and this permission notice shall be included in all
-- copies or substantial portions of the Software.

-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
-- IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
-- FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
-- AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
-- LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
-- OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
-- SOFTWARE.

LIBRARY IEEE; 
USE IEEE.STD_LOGIC_1164.ALL; 
USE IEEE.NUMERIC_STD.ALL; 
  
ENTITY connector IS 
	GENERIC(d : INTEGER := 1000; ----dimentionsize 
	p: INTEGER:= 1000 ); --- prunsize 
	PORT ( 
		input         : IN  STD_LOGIC_VECTOR (d-1 DOWNTO 0); 
		pruneoutput        : OUT  STD_LOGIC_VECTOR (p-1 DOWNTO 0)      
	);
END ENTITY connector;

ARCHITECTURE behavioral OF connector  IS
BEGIN
	 pruneoutput(364) <= input(999);
	 pruneoutput(363) <= input(995);
	 pruneoutput(362) <= input(992);
	 pruneoutput(361) <= input(991);
	 pruneoutput(360) <= input(990);
	 pruneoutput(359) <= input(989);
	 pruneoutput(358) <= input(980);
	 pruneoutput(357) <= input(979);
	 pruneoutput(356) <= input(978);
	 pruneoutput(355) <= input(973);
	 pruneoutput(354) <= input(969);
	 pruneoutput(353) <= input(968);
	 pruneoutput(352) <= input(964);
	 pruneoutput(351) <= input(963);
	 pruneoutput(350) <= input(962);
	 pruneoutput(349) <= input(961);
	 pruneoutput(348) <= input(960);
	 pruneoutput(347) <= input(959);
	 pruneoutput(346) <= input(958);
	 pruneoutput(345) <= input(954);
	 pruneoutput(344) <= input(951);
	 pruneoutput(343) <= input(950);
	 pruneoutput(342) <= input(942);
	 pruneoutput(341) <= input(941);
	 pruneoutput(340) <= input(939);
	 pruneoutput(339) <= input(936);
	 pruneoutput(338) <= input(932);
	 pruneoutput(337) <= input(930);
	 pruneoutput(336) <= input(929);
	 pruneoutput(335) <= input(928);
	 pruneoutput(334) <= input(922);
	 pruneoutput(333) <= input(921);
	 pruneoutput(332) <= input(918);
	 pruneoutput(331) <= input(917);
	 pruneoutput(330) <= input(916);
	 pruneoutput(329) <= input(915);
	 pruneoutput(328) <= input(913);
	 pruneoutput(327) <= input(912);
	 pruneoutput(326) <= input(909);
	 pruneoutput(325) <= input(908);
	 pruneoutput(324) <= input(902);
	 pruneoutput(323) <= input(901);
	 pruneoutput(322) <= input(899);
	 pruneoutput(321) <= input(894);
	 pruneoutput(320) <= input(893);
	 pruneoutput(319) <= input(892);
	 pruneoutput(318) <= input(891);
	 pruneoutput(317) <= input(881);
	 pruneoutput(316) <= input(878);
	 pruneoutput(315) <= input(877);
	 pruneoutput(314) <= input(873);
	 pruneoutput(313) <= input(872);
	 pruneoutput(312) <= input(871);
	 pruneoutput(311) <= input(867);
	 pruneoutput(310) <= input(866);
	 pruneoutput(309) <= input(865);
	 pruneoutput(308) <= input(863);
	 pruneoutput(307) <= input(861);
	 pruneoutput(306) <= input(860);
	 pruneoutput(305) <= input(859);
	 pruneoutput(304) <= input(841);
	 pruneoutput(303) <= input(834);
	 pruneoutput(302) <= input(832);
	 pruneoutput(301) <= input(831);
	 pruneoutput(300) <= input(830);
	 pruneoutput(299) <= input(826);
	 pruneoutput(298) <= input(823);
	 pruneoutput(297) <= input(822);
	 pruneoutput(296) <= input(815);
	 pruneoutput(295) <= input(814);
	 pruneoutput(294) <= input(813);
	 pruneoutput(293) <= input(809);
	 pruneoutput(292) <= input(808);
	 pruneoutput(291) <= input(807);
	 pruneoutput(290) <= input(806);
	 pruneoutput(289) <= input(792);
	 pruneoutput(288) <= input(791);
	 pruneoutput(287) <= input(787);
	 pruneoutput(286) <= input(783);
	 pruneoutput(285) <= input(780);
	 pruneoutput(284) <= input(779);
	 pruneoutput(283) <= input(778);
	 pruneoutput(282) <= input(777);
	 pruneoutput(281) <= input(776);
	 pruneoutput(280) <= input(775);
	 pruneoutput(279) <= input(774);
	 pruneoutput(278) <= input(773);
	 pruneoutput(277) <= input(772);
	 pruneoutput(276) <= input(771);
	 pruneoutput(275) <= input(770);
	 pruneoutput(274) <= input(759);
	 pruneoutput(273) <= input(758);
	 pruneoutput(272) <= input(757);
	 pruneoutput(271) <= input(740);
	 pruneoutput(270) <= input(739);
	 pruneoutput(269) <= input(734);
	 pruneoutput(268) <= input(733);
	 pruneoutput(267) <= input(723);
	 pruneoutput(266) <= input(722);
	 pruneoutput(265) <= input(721);
	 pruneoutput(264) <= input(720);
	 pruneoutput(263) <= input(717);
	 pruneoutput(262) <= input(716);
	 pruneoutput(261) <= input(715);
	 pruneoutput(260) <= input(714);
	 pruneoutput(259) <= input(713);
	 pruneoutput(258) <= input(712);
	 pruneoutput(257) <= input(711);
	 pruneoutput(256) <= input(710);
	 pruneoutput(255) <= input(709);
	 pruneoutput(254) <= input(701);
	 pruneoutput(253) <= input(700);
	 pruneoutput(252) <= input(699);
	 pruneoutput(251) <= input(698);
	 pruneoutput(250) <= input(697);
	 pruneoutput(249) <= input(696);
	 pruneoutput(248) <= input(688);
	 pruneoutput(247) <= input(680);
	 pruneoutput(246) <= input(678);
	 pruneoutput(245) <= input(677);
	 pruneoutput(244) <= input(676);
	 pruneoutput(243) <= input(675);
	 pruneoutput(242) <= input(674);
	 pruneoutput(241) <= input(673);
	 pruneoutput(240) <= input(672);
	 pruneoutput(239) <= input(669);
	 pruneoutput(238) <= input(668);
	 pruneoutput(237) <= input(666);
	 pruneoutput(236) <= input(665);
	 pruneoutput(235) <= input(664);
	 pruneoutput(234) <= input(661);
	 pruneoutput(233) <= input(660);
	 pruneoutput(232) <= input(659);
	 pruneoutput(231) <= input(658);
	 pruneoutput(230) <= input(657);
	 pruneoutput(229) <= input(651);
	 pruneoutput(228) <= input(650);
	 pruneoutput(227) <= input(643);
	 pruneoutput(226) <= input(633);
	 pruneoutput(225) <= input(632);
	 pruneoutput(224) <= input(631);
	 pruneoutput(223) <= input(630);
	 pruneoutput(222) <= input(629);
	 pruneoutput(221) <= input(627);
	 pruneoutput(220) <= input(622);
	 pruneoutput(219) <= input(619);
	 pruneoutput(218) <= input(618);
	 pruneoutput(217) <= input(617);
	 pruneoutput(216) <= input(616);
	 pruneoutput(215) <= input(615);
	 pruneoutput(214) <= input(614);
	 pruneoutput(213) <= input(612);
	 pruneoutput(212) <= input(611);
	 pruneoutput(211) <= input(608);
	 pruneoutput(210) <= input(606);
	 pruneoutput(209) <= input(605);
	 pruneoutput(208) <= input(604);
	 pruneoutput(207) <= input(602);
	 pruneoutput(206) <= input(601);
	 pruneoutput(205) <= input(592);
	 pruneoutput(204) <= input(591);
	 pruneoutput(203) <= input(587);
	 pruneoutput(202) <= input(586);
	 pruneoutput(201) <= input(578);
	 pruneoutput(200) <= input(577);
	 pruneoutput(199) <= input(576);
	 pruneoutput(198) <= input(570);
	 pruneoutput(197) <= input(569);
	 pruneoutput(196) <= input(568);
	 pruneoutput(195) <= input(562);
	 pruneoutput(194) <= input(550);
	 pruneoutput(193) <= input(549);
	 pruneoutput(192) <= input(548);
	 pruneoutput(191) <= input(543);
	 pruneoutput(190) <= input(542);
	 pruneoutput(189) <= input(541);
	 pruneoutput(188) <= input(540);
	 pruneoutput(187) <= input(539);
	 pruneoutput(186) <= input(535);
	 pruneoutput(185) <= input(534);
	 pruneoutput(184) <= input(521);
	 pruneoutput(183) <= input(520);
	 pruneoutput(182) <= input(519);
	 pruneoutput(181) <= input(518);
	 pruneoutput(180) <= input(517);
	 pruneoutput(179) <= input(516);
	 pruneoutput(178) <= input(515);
	 pruneoutput(177) <= input(512);
	 pruneoutput(176) <= input(502);
	 pruneoutput(175) <= input(500);
	 pruneoutput(174) <= input(498);
	 pruneoutput(173) <= input(482);
	 pruneoutput(172) <= input(481);
	 pruneoutput(171) <= input(480);
	 pruneoutput(170) <= input(477);
	 pruneoutput(169) <= input(475);
	 pruneoutput(168) <= input(474);
	 pruneoutput(167) <= input(473);
	 pruneoutput(166) <= input(464);
	 pruneoutput(165) <= input(446);
	 pruneoutput(164) <= input(445);
	 pruneoutput(163) <= input(435);
	 pruneoutput(162) <= input(432);
	 pruneoutput(161) <= input(412);
	 pruneoutput(160) <= input(411);
	 pruneoutput(159) <= input(410);
	 pruneoutput(158) <= input(409);
	 pruneoutput(157) <= input(408);
	 pruneoutput(156) <= input(403);
	 pruneoutput(155) <= input(402);
	 pruneoutput(154) <= input(401);
	 pruneoutput(153) <= input(400);
	 pruneoutput(152) <= input(399);
	 pruneoutput(151) <= input(398);
	 pruneoutput(150) <= input(397);
	 pruneoutput(149) <= input(396);
	 pruneoutput(148) <= input(395);
	 pruneoutput(147) <= input(392);
	 pruneoutput(146) <= input(391);
	 pruneoutput(145) <= input(390);
	 pruneoutput(144) <= input(388);
	 pruneoutput(143) <= input(387);
	 pruneoutput(142) <= input(380);
	 pruneoutput(141) <= input(379);
	 pruneoutput(140) <= input(375);
	 pruneoutput(139) <= input(374);
	 pruneoutput(138) <= input(373);
	 pruneoutput(137) <= input(372);
	 pruneoutput(136) <= input(371);
	 pruneoutput(135) <= input(370);
	 pruneoutput(134) <= input(367);
	 pruneoutput(133) <= input(362);
	 pruneoutput(132) <= input(361);
	 pruneoutput(131) <= input(360);
	 pruneoutput(130) <= input(359);
	 pruneoutput(129) <= input(358);
	 pruneoutput(128) <= input(354);
	 pruneoutput(127) <= input(353);
	 pruneoutput(126) <= input(352);
	 pruneoutput(125) <= input(348);
	 pruneoutput(124) <= input(347);
	 pruneoutput(123) <= input(339);
	 pruneoutput(122) <= input(338);
	 pruneoutput(121) <= input(337);
	 pruneoutput(120) <= input(331);
	 pruneoutput(119) <= input(330);
	 pruneoutput(118) <= input(320);
	 pruneoutput(117) <= input(317);
	 pruneoutput(116) <= input(316);
	 pruneoutput(115) <= input(315);
	 pruneoutput(114) <= input(312);
	 pruneoutput(113) <= input(311);
	 pruneoutput(112) <= input(310);
	 pruneoutput(111) <= input(304);
	 pruneoutput(110) <= input(303);
	 pruneoutput(109) <= input(300);
	 pruneoutput(108) <= input(298);
	 pruneoutput(107) <= input(297);
	 pruneoutput(106) <= input(294);
	 pruneoutput(105) <= input(289);
	 pruneoutput(104) <= input(288);
	 pruneoutput(103) <= input(282);
	 pruneoutput(102) <= input(273);
	 pruneoutput(101) <= input(272);
	 pruneoutput(100) <= input(271);
	 pruneoutput(99) <= input(269);
	 pruneoutput(98) <= input(265);
	 pruneoutput(97) <= input(264);
	 pruneoutput(96) <= input(263);
	 pruneoutput(95) <= input(262);
	 pruneoutput(94) <= input(261);
	 pruneoutput(93) <= input(260);
	 pruneoutput(92) <= input(259);
	 pruneoutput(91) <= input(258);
	 pruneoutput(90) <= input(257);
	 pruneoutput(89) <= input(244);
	 pruneoutput(88) <= input(235);
	 pruneoutput(87) <= input(234);
	 pruneoutput(86) <= input(233);
	 pruneoutput(85) <= input(232);
	 pruneoutput(84) <= input(227);
	 pruneoutput(83) <= input(225);
	 pruneoutput(82) <= input(224);
	 pruneoutput(81) <= input(223);
	 pruneoutput(80) <= input(222);
	 pruneoutput(79) <= input(217);
	 pruneoutput(78) <= input(215);
	 pruneoutput(77) <= input(211);
	 pruneoutput(76) <= input(208);
	 pruneoutput(75) <= input(206);
	 pruneoutput(74) <= input(205);
	 pruneoutput(73) <= input(202);
	 pruneoutput(72) <= input(201);
	 pruneoutput(71) <= input(200);
	 pruneoutput(70) <= input(199);
	 pruneoutput(69) <= input(195);
	 pruneoutput(68) <= input(194);
	 pruneoutput(67) <= input(192);
	 pruneoutput(66) <= input(188);
	 pruneoutput(65) <= input(187);
	 pruneoutput(64) <= input(181);
	 pruneoutput(63) <= input(173);
	 pruneoutput(62) <= input(168);
	 pruneoutput(61) <= input(167);
	 pruneoutput(60) <= input(166);
	 pruneoutput(59) <= input(165);
	 pruneoutput(58) <= input(161);
	 pruneoutput(57) <= input(160);
	 pruneoutput(56) <= input(159);
	 pruneoutput(55) <= input(158);
	 pruneoutput(54) <= input(151);
	 pruneoutput(53) <= input(138);
	 pruneoutput(52) <= input(134);
	 pruneoutput(51) <= input(132);
	 pruneoutput(50) <= input(131);
	 pruneoutput(49) <= input(122);
	 pruneoutput(48) <= input(121);
	 pruneoutput(47) <= input(120);
	 pruneoutput(46) <= input(100);
	 pruneoutput(45) <= input(99);
	 pruneoutput(44) <= input(98);
	 pruneoutput(43) <= input(97);
	 pruneoutput(42) <= input(96);
	 pruneoutput(41) <= input(89);
	 pruneoutput(40) <= input(88);
	 pruneoutput(39) <= input(87);
	 pruneoutput(38) <= input(86);
	 pruneoutput(37) <= input(85);
	 pruneoutput(36) <= input(84);
	 pruneoutput(35) <= input(82);
	 pruneoutput(34) <= input(81);
	 pruneoutput(33) <= input(80);
	 pruneoutput(32) <= input(79);
	 pruneoutput(31) <= input(78);
	 pruneoutput(30) <= input(77);
	 pruneoutput(29) <= input(76);
	 pruneoutput(28) <= input(75);
	 pruneoutput(27) <= input(71);
	 pruneoutput(26) <= input(70);
	 pruneoutput(25) <= input(69);
	 pruneoutput(24) <= input(67);
	 pruneoutput(23) <= input(66);
	 pruneoutput(22) <= input(61);
	 pruneoutput(21) <= input(60);
	 pruneoutput(20) <= input(59);
	 pruneoutput(19) <= input(58);
	 pruneoutput(18) <= input(55);
	 pruneoutput(17) <= input(54);
	 pruneoutput(16) <= input(53);
	 pruneoutput(15) <= input(44);
	 pruneoutput(14) <= input(43);
	 pruneoutput(13) <= input(42);
	 pruneoutput(12) <= input(41);
	 pruneoutput(11) <= input(31);
	 pruneoutput(10) <= input(30);
	 pruneoutput(9) <= input(29);
	 pruneoutput(8) <= input(28);
	 pruneoutput(7) <= input(23);
	 pruneoutput(6) <= input(16);
	 pruneoutput(5) <= input(15);
	 pruneoutput(4) <= input(14);
	 pruneoutput(3) <= input(9);
	 pruneoutput(2) <= input(5);
	 pruneoutput(1) <= input(1);
	 pruneoutput(0) <= input(0);

END ARCHITECTURE behavioral;