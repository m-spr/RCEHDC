LIBRARY IEEE; 
USE IEEE.STD_LOGIC_1164.ALL; 
USE IEEE.NUMERIC_STD.ALL; 
  
ENTITY connector IS 
	PORT ( 
		input         : IN  STD_LOGIC_VECTOR (999 DOWNTO 0); 
		pruneoutput        : OUT  STD_LOGIC_VECTOR (665 DOWNTO 0)      
	);
END ENTITY connector;

ARCHITECTURE behavioral OF connector  IS
BEGIN
pruneoutput(0) <= input(0);
pruneoutput(1) <= input(5);
pruneoutput(2) <= input(7);
pruneoutput(3) <= input(8);
pruneoutput(4) <= input(10);
pruneoutput(5) <= input(16);
pruneoutput(6) <= input(19);
pruneoutput(7) <= input(24);
pruneoutput(8) <= input(25);
pruneoutput(9) <= input(26);
pruneoutput(10) <= input(31);
pruneoutput(11) <= input(38);
pruneoutput(12) <= input(39);
pruneoutput(13) <= input(40);
pruneoutput(14) <= input(41);
pruneoutput(15) <= input(42);
pruneoutput(16) <= input(46);
pruneoutput(17) <= input(48);
pruneoutput(18) <= input(49);
pruneoutput(19) <= input(50);
pruneoutput(20) <= input(52);
pruneoutput(21) <= input(53);
pruneoutput(22) <= input(54);
pruneoutput(23) <= input(57);
pruneoutput(24) <= input(58);
pruneoutput(25) <= input(59);
pruneoutput(26) <= input(60);
pruneoutput(27) <= input(61);
pruneoutput(28) <= input(63);
pruneoutput(29) <= input(64);
pruneoutput(30) <= input(69);
pruneoutput(31) <= input(70);
pruneoutput(32) <= input(71);
pruneoutput(33) <= input(72);
pruneoutput(34) <= input(74);
pruneoutput(35) <= input(75);
pruneoutput(36) <= input(76);
pruneoutput(37) <= input(77);
pruneoutput(38) <= input(79);
pruneoutput(39) <= input(80);
pruneoutput(40) <= input(81);
pruneoutput(41) <= input(82);
pruneoutput(42) <= input(83);
pruneoutput(43) <= input(84);
pruneoutput(44) <= input(85);
pruneoutput(45) <= input(86);
pruneoutput(46) <= input(87);
pruneoutput(47) <= input(88);
pruneoutput(48) <= input(90);
pruneoutput(49) <= input(91);
pruneoutput(50) <= input(93);
pruneoutput(51) <= input(94);
pruneoutput(52) <= input(95);
pruneoutput(53) <= input(96);
pruneoutput(54) <= input(97);
pruneoutput(55) <= input(98);
pruneoutput(56) <= input(99);
pruneoutput(57) <= input(103);
pruneoutput(58) <= input(104);
pruneoutput(59) <= input(108);
pruneoutput(60) <= input(109);
pruneoutput(61) <= input(110);
pruneoutput(62) <= input(111);
pruneoutput(63) <= input(112);
pruneoutput(64) <= input(113);
pruneoutput(65) <= input(114);
pruneoutput(66) <= input(115);
pruneoutput(67) <= input(116);
pruneoutput(68) <= input(117);
pruneoutput(69) <= input(118);
pruneoutput(70) <= input(119);
pruneoutput(71) <= input(120);
pruneoutput(72) <= input(121);
pruneoutput(73) <= input(126);
pruneoutput(74) <= input(128);
pruneoutput(75) <= input(129);
pruneoutput(76) <= input(130);
pruneoutput(77) <= input(131);
pruneoutput(78) <= input(132);
pruneoutput(79) <= input(133);
pruneoutput(80) <= input(134);
pruneoutput(81) <= input(136);
pruneoutput(82) <= input(137);
pruneoutput(83) <= input(138);
pruneoutput(84) <= input(139);
pruneoutput(85) <= input(141);
pruneoutput(86) <= input(142);
pruneoutput(87) <= input(143);
pruneoutput(88) <= input(144);
pruneoutput(89) <= input(145);
pruneoutput(90) <= input(146);
pruneoutput(91) <= input(147);
pruneoutput(92) <= input(148);
pruneoutput(93) <= input(149);
pruneoutput(94) <= input(150);
pruneoutput(95) <= input(151);
pruneoutput(96) <= input(152);
pruneoutput(97) <= input(153);
pruneoutput(98) <= input(154);
pruneoutput(99) <= input(155);
pruneoutput(100) <= input(157);
pruneoutput(101) <= input(158);
pruneoutput(102) <= input(159);
pruneoutput(103) <= input(160);
pruneoutput(104) <= input(161);
pruneoutput(105) <= input(162);
pruneoutput(106) <= input(165);
pruneoutput(107) <= input(166);
pruneoutput(108) <= input(168);
pruneoutput(109) <= input(170);
pruneoutput(110) <= input(171);
pruneoutput(111) <= input(172);
pruneoutput(112) <= input(173);
pruneoutput(113) <= input(174);
pruneoutput(114) <= input(175);
pruneoutput(115) <= input(178);
pruneoutput(116) <= input(179);
pruneoutput(117) <= input(182);
pruneoutput(118) <= input(183);
pruneoutput(119) <= input(184);
pruneoutput(120) <= input(185);
pruneoutput(121) <= input(186);
pruneoutput(122) <= input(188);
pruneoutput(123) <= input(189);
pruneoutput(124) <= input(190);
pruneoutput(125) <= input(191);
pruneoutput(126) <= input(192);
pruneoutput(127) <= input(193);
pruneoutput(128) <= input(194);
pruneoutput(129) <= input(197);
pruneoutput(130) <= input(198);
pruneoutput(131) <= input(199);
pruneoutput(132) <= input(200);
pruneoutput(133) <= input(205);
pruneoutput(134) <= input(209);
pruneoutput(135) <= input(210);
pruneoutput(136) <= input(212);
pruneoutput(137) <= input(213);
pruneoutput(138) <= input(216);
pruneoutput(139) <= input(217);
pruneoutput(140) <= input(220);
pruneoutput(141) <= input(221);
pruneoutput(142) <= input(222);
pruneoutput(143) <= input(225);
pruneoutput(144) <= input(226);
pruneoutput(145) <= input(231);
pruneoutput(146) <= input(232);
pruneoutput(147) <= input(235);
pruneoutput(148) <= input(236);
pruneoutput(149) <= input(237);
pruneoutput(150) <= input(240);
pruneoutput(151) <= input(241);
pruneoutput(152) <= input(242);
pruneoutput(153) <= input(245);
pruneoutput(154) <= input(246);
pruneoutput(155) <= input(248);
pruneoutput(156) <= input(253);
pruneoutput(157) <= input(255);
pruneoutput(158) <= input(256);
pruneoutput(159) <= input(257);
pruneoutput(160) <= input(258);
pruneoutput(161) <= input(264);
pruneoutput(162) <= input(265);
pruneoutput(163) <= input(266);
pruneoutput(164) <= input(267);
pruneoutput(165) <= input(269);
pruneoutput(166) <= input(270);
pruneoutput(167) <= input(271);
pruneoutput(168) <= input(272);
pruneoutput(169) <= input(273);
pruneoutput(170) <= input(274);
pruneoutput(171) <= input(275);
pruneoutput(172) <= input(276);
pruneoutput(173) <= input(278);
pruneoutput(174) <= input(279);
pruneoutput(175) <= input(281);
pruneoutput(176) <= input(285);
pruneoutput(177) <= input(286);
pruneoutput(178) <= input(287);
pruneoutput(179) <= input(288);
pruneoutput(180) <= input(289);
pruneoutput(181) <= input(290);
pruneoutput(182) <= input(291);
pruneoutput(183) <= input(296);
pruneoutput(184) <= input(299);
pruneoutput(185) <= input(301);
pruneoutput(186) <= input(302);
pruneoutput(187) <= input(303);
pruneoutput(188) <= input(304);
pruneoutput(189) <= input(305);
pruneoutput(190) <= input(306);
pruneoutput(191) <= input(307);
pruneoutput(192) <= input(308);
pruneoutput(193) <= input(310);
pruneoutput(194) <= input(312);
pruneoutput(195) <= input(313);
pruneoutput(196) <= input(314);
pruneoutput(197) <= input(315);
pruneoutput(198) <= input(316);
pruneoutput(199) <= input(317);
pruneoutput(200) <= input(318);
pruneoutput(201) <= input(319);
pruneoutput(202) <= input(320);
pruneoutput(203) <= input(321);
pruneoutput(204) <= input(322);
pruneoutput(205) <= input(323);
pruneoutput(206) <= input(328);
pruneoutput(207) <= input(334);
pruneoutput(208) <= input(335);
pruneoutput(209) <= input(336);
pruneoutput(210) <= input(337);
pruneoutput(211) <= input(338);
pruneoutput(212) <= input(339);
pruneoutput(213) <= input(340);
pruneoutput(214) <= input(342);
pruneoutput(215) <= input(343);
pruneoutput(216) <= input(346);
pruneoutput(217) <= input(347);
pruneoutput(218) <= input(348);
pruneoutput(219) <= input(349);
pruneoutput(220) <= input(355);
pruneoutput(221) <= input(356);
pruneoutput(222) <= input(357);
pruneoutput(223) <= input(358);
pruneoutput(224) <= input(359);
pruneoutput(225) <= input(360);
pruneoutput(226) <= input(361);
pruneoutput(227) <= input(362);
pruneoutput(228) <= input(363);
pruneoutput(229) <= input(364);
pruneoutput(230) <= input(366);
pruneoutput(231) <= input(367);
pruneoutput(232) <= input(368);
pruneoutput(233) <= input(369);
pruneoutput(234) <= input(370);
pruneoutput(235) <= input(371);
pruneoutput(236) <= input(372);
pruneoutput(237) <= input(377);
pruneoutput(238) <= input(378);
pruneoutput(239) <= input(379);
pruneoutput(240) <= input(380);
pruneoutput(241) <= input(381);
pruneoutput(242) <= input(382);
pruneoutput(243) <= input(384);
pruneoutput(244) <= input(387);
pruneoutput(245) <= input(388);
pruneoutput(246) <= input(393);
pruneoutput(247) <= input(394);
pruneoutput(248) <= input(395);
pruneoutput(249) <= input(396);
pruneoutput(250) <= input(397);
pruneoutput(251) <= input(398);
pruneoutput(252) <= input(399);
pruneoutput(253) <= input(400);
pruneoutput(254) <= input(401);
pruneoutput(255) <= input(402);
pruneoutput(256) <= input(403);
pruneoutput(257) <= input(404);
pruneoutput(258) <= input(405);
pruneoutput(259) <= input(406);
pruneoutput(260) <= input(412);
pruneoutput(261) <= input(413);
pruneoutput(262) <= input(414);
pruneoutput(263) <= input(417);
pruneoutput(264) <= input(418);
pruneoutput(265) <= input(419);
pruneoutput(266) <= input(420);
pruneoutput(267) <= input(421);
pruneoutput(268) <= input(422);
pruneoutput(269) <= input(423);
pruneoutput(270) <= input(425);
pruneoutput(271) <= input(426);
pruneoutput(272) <= input(427);
pruneoutput(273) <= input(428);
pruneoutput(274) <= input(429);
pruneoutput(275) <= input(430);
pruneoutput(276) <= input(431);
pruneoutput(277) <= input(432);
pruneoutput(278) <= input(433);
pruneoutput(279) <= input(434);
pruneoutput(280) <= input(435);
pruneoutput(281) <= input(436);
pruneoutput(282) <= input(437);
pruneoutput(283) <= input(438);
pruneoutput(284) <= input(439);
pruneoutput(285) <= input(440);
pruneoutput(286) <= input(441);
pruneoutput(287) <= input(442);
pruneoutput(288) <= input(443);
pruneoutput(289) <= input(444);
pruneoutput(290) <= input(445);
pruneoutput(291) <= input(446);
pruneoutput(292) <= input(447);
pruneoutput(293) <= input(448);
pruneoutput(294) <= input(450);
pruneoutput(295) <= input(451);
pruneoutput(296) <= input(452);
pruneoutput(297) <= input(453);
pruneoutput(298) <= input(454);
pruneoutput(299) <= input(455);
pruneoutput(300) <= input(456);
pruneoutput(301) <= input(462);
pruneoutput(302) <= input(463);
pruneoutput(303) <= input(466);
pruneoutput(304) <= input(470);
pruneoutput(305) <= input(478);
pruneoutput(306) <= input(480);
pruneoutput(307) <= input(484);
pruneoutput(308) <= input(485);
pruneoutput(309) <= input(486);
pruneoutput(310) <= input(487);
pruneoutput(311) <= input(488);
pruneoutput(312) <= input(489);
pruneoutput(313) <= input(490);
pruneoutput(314) <= input(491);
pruneoutput(315) <= input(492);
pruneoutput(316) <= input(493);
pruneoutput(317) <= input(494);
pruneoutput(318) <= input(498);
pruneoutput(319) <= input(500);
pruneoutput(320) <= input(501);
pruneoutput(321) <= input(503);
pruneoutput(322) <= input(504);
pruneoutput(323) <= input(505);
pruneoutput(324) <= input(506);
pruneoutput(325) <= input(507);
pruneoutput(326) <= input(508);
pruneoutput(327) <= input(509);
pruneoutput(328) <= input(515);
pruneoutput(329) <= input(516);
pruneoutput(330) <= input(517);
pruneoutput(331) <= input(518);
pruneoutput(332) <= input(519);
pruneoutput(333) <= input(520);
pruneoutput(334) <= input(524);
pruneoutput(335) <= input(525);
pruneoutput(336) <= input(526);
pruneoutput(337) <= input(527);
pruneoutput(338) <= input(528);
pruneoutput(339) <= input(529);
pruneoutput(340) <= input(530);
pruneoutput(341) <= input(531);
pruneoutput(342) <= input(532);
pruneoutput(343) <= input(540);
pruneoutput(344) <= input(541);
pruneoutput(345) <= input(544);
pruneoutput(346) <= input(545);
pruneoutput(347) <= input(547);
pruneoutput(348) <= input(549);
pruneoutput(349) <= input(550);
pruneoutput(350) <= input(557);
pruneoutput(351) <= input(558);
pruneoutput(352) <= input(559);
pruneoutput(353) <= input(560);
pruneoutput(354) <= input(561);
pruneoutput(355) <= input(562);
pruneoutput(356) <= input(563);
pruneoutput(357) <= input(564);
pruneoutput(358) <= input(565);
pruneoutput(359) <= input(566);
pruneoutput(360) <= input(567);
pruneoutput(361) <= input(568);
pruneoutput(362) <= input(569);
pruneoutput(363) <= input(570);
pruneoutput(364) <= input(571);
pruneoutput(365) <= input(572);
pruneoutput(366) <= input(573);
pruneoutput(367) <= input(574);
pruneoutput(368) <= input(575);
pruneoutput(369) <= input(576);
pruneoutput(370) <= input(581);
pruneoutput(371) <= input(582);
pruneoutput(372) <= input(583);
pruneoutput(373) <= input(584);
pruneoutput(374) <= input(585);
pruneoutput(375) <= input(588);
pruneoutput(376) <= input(590);
pruneoutput(377) <= input(594);
pruneoutput(378) <= input(595);
pruneoutput(379) <= input(596);
pruneoutput(380) <= input(598);
pruneoutput(381) <= input(599);
pruneoutput(382) <= input(601);
pruneoutput(383) <= input(602);
pruneoutput(384) <= input(603);
pruneoutput(385) <= input(608);
pruneoutput(386) <= input(609);
pruneoutput(387) <= input(610);
pruneoutput(388) <= input(611);
pruneoutput(389) <= input(612);
pruneoutput(390) <= input(613);
pruneoutput(391) <= input(614);
pruneoutput(392) <= input(615);
pruneoutput(393) <= input(616);
pruneoutput(394) <= input(617);
pruneoutput(395) <= input(618);
pruneoutput(396) <= input(621);
pruneoutput(397) <= input(624);
pruneoutput(398) <= input(625);
pruneoutput(399) <= input(626);
pruneoutput(400) <= input(627);
pruneoutput(401) <= input(629);
pruneoutput(402) <= input(630);
pruneoutput(403) <= input(631);
pruneoutput(404) <= input(632);
pruneoutput(405) <= input(633);
pruneoutput(406) <= input(634);
pruneoutput(407) <= input(635);
pruneoutput(408) <= input(636);
pruneoutput(409) <= input(637);
pruneoutput(410) <= input(638);
pruneoutput(411) <= input(639);
pruneoutput(412) <= input(640);
pruneoutput(413) <= input(641);
pruneoutput(414) <= input(642);
pruneoutput(415) <= input(643);
pruneoutput(416) <= input(644);
pruneoutput(417) <= input(645);
pruneoutput(418) <= input(646);
pruneoutput(419) <= input(647);
pruneoutput(420) <= input(648);
pruneoutput(421) <= input(649);
pruneoutput(422) <= input(650);
pruneoutput(423) <= input(651);
pruneoutput(424) <= input(655);
pruneoutput(425) <= input(656);
pruneoutput(426) <= input(660);
pruneoutput(427) <= input(661);
pruneoutput(428) <= input(663);
pruneoutput(429) <= input(664);
pruneoutput(430) <= input(665);
pruneoutput(431) <= input(666);
pruneoutput(432) <= input(667);
pruneoutput(433) <= input(668);
pruneoutput(434) <= input(669);
pruneoutput(435) <= input(672);
pruneoutput(436) <= input(673);
pruneoutput(437) <= input(674);
pruneoutput(438) <= input(675);
pruneoutput(439) <= input(676);
pruneoutput(440) <= input(677);
pruneoutput(441) <= input(678);
pruneoutput(442) <= input(679);
pruneoutput(443) <= input(680);
pruneoutput(444) <= input(681);
pruneoutput(445) <= input(685);
pruneoutput(446) <= input(686);
pruneoutput(447) <= input(687);
pruneoutput(448) <= input(688);
pruneoutput(449) <= input(693);
pruneoutput(450) <= input(694);
pruneoutput(451) <= input(695);
pruneoutput(452) <= input(696);
pruneoutput(453) <= input(705);
pruneoutput(454) <= input(710);
pruneoutput(455) <= input(711);
pruneoutput(456) <= input(712);
pruneoutput(457) <= input(714);
pruneoutput(458) <= input(720);
pruneoutput(459) <= input(721);
pruneoutput(460) <= input(723);
pruneoutput(461) <= input(730);
pruneoutput(462) <= input(734);
pruneoutput(463) <= input(735);
pruneoutput(464) <= input(736);
pruneoutput(465) <= input(737);
pruneoutput(466) <= input(738);
pruneoutput(467) <= input(739);
pruneoutput(468) <= input(740);
pruneoutput(469) <= input(745);
pruneoutput(470) <= input(749);
pruneoutput(471) <= input(750);
pruneoutput(472) <= input(751);
pruneoutput(473) <= input(752);
pruneoutput(474) <= input(753);
pruneoutput(475) <= input(754);
pruneoutput(476) <= input(755);
pruneoutput(477) <= input(758);
pruneoutput(478) <= input(759);
pruneoutput(479) <= input(760);
pruneoutput(480) <= input(761);
pruneoutput(481) <= input(762);
pruneoutput(482) <= input(763);
pruneoutput(483) <= input(764);
pruneoutput(484) <= input(766);
pruneoutput(485) <= input(767);
pruneoutput(486) <= input(768);
pruneoutput(487) <= input(769);
pruneoutput(488) <= input(770);
pruneoutput(489) <= input(774);
pruneoutput(490) <= input(776);
pruneoutput(491) <= input(777);
pruneoutput(492) <= input(778);
pruneoutput(493) <= input(780);
pruneoutput(494) <= input(781);
pruneoutput(495) <= input(782);
pruneoutput(496) <= input(783);
pruneoutput(497) <= input(784);
pruneoutput(498) <= input(785);
pruneoutput(499) <= input(792);
pruneoutput(500) <= input(793);
pruneoutput(501) <= input(794);
pruneoutput(502) <= input(796);
pruneoutput(503) <= input(798);
pruneoutput(504) <= input(799);
pruneoutput(505) <= input(800);
pruneoutput(506) <= input(802);
pruneoutput(507) <= input(803);
pruneoutput(508) <= input(804);
pruneoutput(509) <= input(805);
pruneoutput(510) <= input(806);
pruneoutput(511) <= input(807);
pruneoutput(512) <= input(808);
pruneoutput(513) <= input(809);
pruneoutput(514) <= input(810);
pruneoutput(515) <= input(811);
pruneoutput(516) <= input(812);
pruneoutput(517) <= input(813);
pruneoutput(518) <= input(814);
pruneoutput(519) <= input(816);
pruneoutput(520) <= input(817);
pruneoutput(521) <= input(818);
pruneoutput(522) <= input(819);
pruneoutput(523) <= input(820);
pruneoutput(524) <= input(821);
pruneoutput(525) <= input(824);
pruneoutput(526) <= input(825);
pruneoutput(527) <= input(826);
pruneoutput(528) <= input(827);
pruneoutput(529) <= input(832);
pruneoutput(530) <= input(833);
pruneoutput(531) <= input(834);
pruneoutput(532) <= input(837);
pruneoutput(533) <= input(838);
pruneoutput(534) <= input(839);
pruneoutput(535) <= input(842);
pruneoutput(536) <= input(843);
pruneoutput(537) <= input(844);
pruneoutput(538) <= input(845);
pruneoutput(539) <= input(846);
pruneoutput(540) <= input(847);
pruneoutput(541) <= input(850);
pruneoutput(542) <= input(851);
pruneoutput(543) <= input(852);
pruneoutput(544) <= input(853);
pruneoutput(545) <= input(854);
pruneoutput(546) <= input(855);
pruneoutput(547) <= input(856);
pruneoutput(548) <= input(857);
pruneoutput(549) <= input(858);
pruneoutput(550) <= input(859);
pruneoutput(551) <= input(860);
pruneoutput(552) <= input(861);
pruneoutput(553) <= input(862);
pruneoutput(554) <= input(863);
pruneoutput(555) <= input(866);
pruneoutput(556) <= input(867);
pruneoutput(557) <= input(869);
pruneoutput(558) <= input(870);
pruneoutput(559) <= input(871);
pruneoutput(560) <= input(874);
pruneoutput(561) <= input(875);
pruneoutput(562) <= input(877);
pruneoutput(563) <= input(878);
pruneoutput(564) <= input(879);
pruneoutput(565) <= input(880);
pruneoutput(566) <= input(881);
pruneoutput(567) <= input(882);
pruneoutput(568) <= input(883);
pruneoutput(569) <= input(884);
pruneoutput(570) <= input(885);
pruneoutput(571) <= input(886);
pruneoutput(572) <= input(887);
pruneoutput(573) <= input(890);
pruneoutput(574) <= input(891);
pruneoutput(575) <= input(892);
pruneoutput(576) <= input(894);
pruneoutput(577) <= input(895);
pruneoutput(578) <= input(896);
pruneoutput(579) <= input(899);
pruneoutput(580) <= input(900);
pruneoutput(581) <= input(901);
pruneoutput(582) <= input(902);
pruneoutput(583) <= input(903);
pruneoutput(584) <= input(904);
pruneoutput(585) <= input(905);
pruneoutput(586) <= input(906);
pruneoutput(587) <= input(907);
pruneoutput(588) <= input(908);
pruneoutput(589) <= input(909);
pruneoutput(590) <= input(910);
pruneoutput(591) <= input(911);
pruneoutput(592) <= input(912);
pruneoutput(593) <= input(913);
pruneoutput(594) <= input(914);
pruneoutput(595) <= input(915);
pruneoutput(596) <= input(916);
pruneoutput(597) <= input(917);
pruneoutput(598) <= input(919);
pruneoutput(599) <= input(920);
pruneoutput(600) <= input(922);
pruneoutput(601) <= input(923);
pruneoutput(602) <= input(924);
pruneoutput(603) <= input(925);
pruneoutput(604) <= input(926);
pruneoutput(605) <= input(932);
pruneoutput(606) <= input(933);
pruneoutput(607) <= input(934);
pruneoutput(608) <= input(935);
pruneoutput(609) <= input(936);
pruneoutput(610) <= input(937);
pruneoutput(611) <= input(938);
pruneoutput(612) <= input(939);
pruneoutput(613) <= input(941);
pruneoutput(614) <= input(942);
pruneoutput(615) <= input(945);
pruneoutput(616) <= input(946);
pruneoutput(617) <= input(947);
pruneoutput(618) <= input(948);
pruneoutput(619) <= input(949);
pruneoutput(620) <= input(950);
pruneoutput(621) <= input(952);
pruneoutput(622) <= input(953);
pruneoutput(623) <= input(954);
pruneoutput(624) <= input(955);
pruneoutput(625) <= input(956);
pruneoutput(626) <= input(957);
pruneoutput(627) <= input(961);
pruneoutput(628) <= input(962);
pruneoutput(629) <= input(963);
pruneoutput(630) <= input(964);
pruneoutput(631) <= input(965);
pruneoutput(632) <= input(966);
pruneoutput(633) <= input(967);
pruneoutput(634) <= input(968);
pruneoutput(635) <= input(969);
pruneoutput(636) <= input(970);
pruneoutput(637) <= input(971);
pruneoutput(638) <= input(972);
pruneoutput(639) <= input(973);
pruneoutput(640) <= input(974);
pruneoutput(641) <= input(975);
pruneoutput(642) <= input(976);
pruneoutput(643) <= input(977);
pruneoutput(644) <= input(978);
pruneoutput(645) <= input(979);
pruneoutput(646) <= input(980);
pruneoutput(647) <= input(981);
pruneoutput(648) <= input(982);
pruneoutput(649) <= input(983);
pruneoutput(650) <= input(984);
pruneoutput(651) <= input(985);
pruneoutput(652) <= input(986);
pruneoutput(653) <= input(987);
pruneoutput(654) <= input(988);
pruneoutput(655) <= input(989);
pruneoutput(656) <= input(990);
pruneoutput(657) <= input(991);
pruneoutput(658) <= input(992);
pruneoutput(659) <= input(993);
pruneoutput(660) <= input(994);
pruneoutput(661) <= input(995);
pruneoutput(662) <= input(996);
pruneoutput(663) <= input(997);
pruneoutput(664) <= input(998);
pruneoutput(665) <= input(999);

END ARCHITECTURE behavioral;