LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY BasedVectorLFSR IS
	GENERIC ( n	: INTEGER	:= 2000			    -- number of bits
				);	 
	PORT (
		clk, rst, update	: IN STD_LOGIC; 
		congigSignitureIn , congigInitialvaluesIn : IN STD_LOGIC_VECTOR (n-1 DOWNTO 0 );
		dout				: OUT  STD_LOGIC_VECTOR (n-1 DOWNTO 0 )
	);
END ENTITY BasedVectorLFSR;

ARCHITECTURE behavioral OF BasedVectorLFSR IS

COMPONENT  regOne IS
	GENERIC (init : STD_LOGIC := '1');   -- initial value
	PORT (
		clk 				: IN  STD_LOGIC;
		regUpdate, regrst 	: IN  STD_LOGIC;
		din        			: IN  STD_LOGIC;
		dout        		: OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL interValIn : STD_LOGIC_VECTOR (n-1 DOWNTO 0);
SIGNAL interValOut : STD_LOGIC_VECTOR (n-1 DOWNTO 0);
SIGNAL interValOutR : STD_LOGIC_VECTOR (0 TO n-1);
CONSTANT congigSigniture : STD_LOGIC_VECTOR (n-1 DOWNTO 0) :=    "1011101110111010011001010011110111001001011001010010110000010101010100001010111001011010010100111111101101011011000110101111010110100000111101011100101011110001110011011001010110001010101100111111010001000000101110001101010100111000010111111111111010001011101101000110101110111100111000010011000110000101011110000001011101010101111000001011011100000110100100110000001000111010100100000000101101000110101110011101111000001011100001000100110000001111011100111111000011001100101011110111001101010010100101011101100011100010111011110001000111001001100010101011100100001000011100011111001110011111001100101111000111110110110001011010101110001110011011110000101100001010001110110000101100110001101001101011111000101011000001100100110101101000111001001001110011111111000101110001100110101001001001000101101110111101100011001010010001101011100010011011010100110100010101110001111011101101000110111010101110101010010001101000111011111101001000000100101101101000001110110000111011100000110111011000111100001110"; --"1010101011000011001011001000001001000110100100000010011011000001110101100010000001000111100011101100011001100110100010101100010001011111010110000011000010111011110110101000110101100100110110100001010010111100101010101000111011111101101111011111001111001010110000010110100001111110011100100000000110110110000000011011010111101011100110101100010100100011010011000001010111000000010001101101101011010110110011110000010000110110010110100011111001011110011010011101011010111100011001010111011111110101100110001110000011111111110110001011001111111110010101010010011101000011100111101011011000110101010101100000100001101010101000111111001001111101010000110001110110001010111000101100101010011110010101100010011011011111111100100111100010011100101010010000001100111011100101101011100010111001000110101111110111111010001000100101100011100010001011001100110111011010101010000010100000000101001000110011011011011100010011011001001011100000000000000001000010010101100101110110001001101010101101010001110000001100";

CONSTANT congigInitialvalues : STD_LOGIC_VECTOR (n-1 DOWNTO 0) := "0110000001110110001111110010001000101100000101110111101011100111101100101100100000011000111100001011110110101111011011001001111010010000011101000110011110110101010001100011111101001100010011000101101110110111101010110111000111101110101100010010001100010010010011010010101111100110110000001011111000100111110011111111110001100111011100011101000110100101100100001001101000001101001111010110010001110101000011100000101101011111101001000101010000100010001100000011001100000001011001001010110111111010011011010000111111101000000101001010111010111000010001111000000110100011101101001100001110010011111000010001001010101100011000101101101100111111100111101011000101110001111011001110110010111101110111010110100100110101001100001100101111000101111101000010100010000010010100100000111110010101010111011011010110101100010010101100100111110111001101000111100101100011100111110011101101000011100010000100011110001100111011001101011100011010010011000001111000101100010110011110000010100001011110111010111011001010";--"1111000000100110110100000110111010000101111100010011000110000110000100100100100010111110100100111000000001010111001001001000111010011010000001011010010100111000100010110111010111110010000101010100011101011111011100001011010100011100110110100001101100111100101111001001100100000011110111000110111000010001111100011110001110001010001011011011000000001010000001000001000011100010110011111101111000000010000111110001101011110111101010101010001110110110100100101011011011011110000111110110011000100110111010000011101100111010000010101011010111001011110110100000101100101111110011010011010010111000100100101100101101010001001110100010100001011100010111110010110011101000111110110001100100011100001110110000101111110011100100011011011101101110010101000101010100101011110011100100111100010011011100100101001010000110000101011100001110011111100011000011101010100001011010100101011110000100010001101001000000001011010001001001001000111010110101000010101011111110000010001010100111111100100011000110110101100110";

BEGIN

	regArr : FOR i IN 1 TO n-1 GENERATE
		Ireg : regOne 
			GENERIC map(congigInitialvalues(i))
			PORT map(clk,  update, rst, 
			interValIn(i), 	interValOut(i) 
					 );   
	END GENERATE regArr;
	xorchain : FOR i IN 1 TO n-1 GENERATE
	xorchain1: IF (congigSigniture(i) = '1') GENERATE
			interValIn(i) <= interValOut(i-1) XOR  interValOut(n-1);
		END GENERATE xorchain1;
	xorchain2: IF (congigSigniture(i) = '0') GENERATE
			interValIn(i) <= interValOut(i-1);
		END GENERATE xorchain2;
	END GENERATE xorchain;
	interValIn(0) <= interValOut(n-1);
	reg0 : regOne 
			GENERIC map(congigInitialvalues(0))
			PORT map(clk,  update, rst, 
			interValIn(0), 	interValOut(0) 
					 ); 
	--interValOutR <= interValOut;
	dout <= interValOut;--(0 TO n-1);

END ARCHITECTURE behavioral;